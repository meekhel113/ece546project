* PEX netlist file	Thu Apr 21 18:10:59 2022	top_level
* icv_netlist Version RHEL64 S-2021.06-SP2.6831572 2021/08/30
*.UNIT=4000

* Hierarchy Level 4
.subckt fill_sram_inverted 2 3 4 5
.ends fill_sram_inverted
.subckt fill_sram 2 3 4 5
.ends fill_sram
.subckt fill_sram_column_decoder_write 2 3 4 5
.ends fill_sram_column_decoder_write
.subckt fill_sram_inverted_read 2 3 4 5
.ends fill_sram_inverted_read
.subckt inverter_row_decoder 2 3 4 5 6 7
.ends inverter_row_decoder
.subckt inverter_column_decoder_write 2 3 4 5 6 7
.ends inverter_column_decoder_write
.subckt sram_6T_1finger_inverted 2 3 4 5 6 7 8 9 10
*.floating_nets _GENERATED_11 _GENERATED_12
.ends sram_6T_1finger_inverted
.subckt sram_6T_1finger 2 3 4 5 6 7 8 9 10
*.floating_nets _GENERATED_11 _GENERATED_12
.ends sram_6T_1finger
.subckt fill_sram_nmos 2 3 4 5 6 7 8
.ends fill_sram_nmos
.subckt inverter_buf_top_leve 2 3 4 5 6 7
.ends inverter_buf_top_leve
.subckt inverter_buf_top_level_v1 2 3 4 5 6 7 8
.ends inverter_buf_top_level_v1
.subckt fill_sram_inverted_pmos_read 2 3 4 5 6
.ends fill_sram_inverted_pmos_read
.subckt fill_sram_pmos 2 3 4 5 6
*.floating_nets _GENERATED_7
.ends fill_sram_pmos
.subckt fill_sram_inverted_nmos 2 3 4 5
.ends fill_sram_inverted_nmos
.subckt and 2 3 4 5 6 7 8 9 10 11
MM1 3 2 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=504 $Y=326  $PIN_XY=(534,508,534,338),504,326,(474,508,474,338) $DEVICE_ID=1003
MM2 6 5 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=336 $Y=326  $PIN_XY=(366,508,366,338),336,326,(306,508,306,338) $DEVICE_ID=1003
MM3 2 4 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=168 $Y=326  $PIN_XY=(198,508,198,338),168,326,(138,508,138,338) $DEVICE_ID=1003
.ends and
.subckt and_v1 2 3 4 5 6 7 8 9 10 11
MM1 3 2 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=504 $Y=326  $PIN_XY=(534,508,534,338),504,326,(474,508,474,338) $DEVICE_ID=1003
MM2 6 5 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=336 $Y=326  $PIN_XY=(366,508,366,338),336,326,(306,508,306,338) $DEVICE_ID=1003
MM3 2 4 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=168 $Y=326  $PIN_XY=(198,508,198,338),168,326,(138,508,138,338) $DEVICE_ID=1003
.ends and_v1
.subckt fill_sram_inverted_pmos_write 2 3 4 5 6
*.floating_nets _GENERATED_7
.ends fill_sram_inverted_pmos_write
.subckt inverter_write 2 3 4 5 6 7 8
MM1 3 2 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=222 $Y=310  $PIN_XY=(252,492,252,322),222,310,(192,492,192,322) $DEVICE_ID=1003
.ends inverter_write
.subckt fill_sram_inverted_write_pmos 2 3 4 5
.ends fill_sram_inverted_write_pmos

* Hierarchy Level 3
.subckt sram_lvs_grid 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 23
+	24 25 26 27 28
XX73A2B172271_1 3 2 4 17 fill_sram_column_decoder_write $T=16 13150 0 0 $X=-8 $Y=13086
XX73A2B172271_2 3 2 4 17 fill_sram_column_decoder_write $T=184 13150 0 0 $X=160 $Y=13086
XX73A2B172273_1 3 2 5 18 fill_sram_inverted $T=16 11840 1 0 $X=-8 $Y=11124
XX73A2B172273_2 3 2 5 18 fill_sram_inverted $T=184 11840 1 0 $X=160 $Y=11124
XX73A2B172275_1 3 2 6 17 fill_sram_inverted $T=16 14456 1 0 $X=-8 $Y=13740
XX73A2B172275_2 3 2 6 17 fill_sram_inverted $T=184 14456 1 0 $X=160 $Y=13740
XX73A2B172277_1 3 2 4 19 fill_sram_inverted $T=16 13148 1 0 $X=-8 $Y=12432
XX73A2B172277_2 3 2 4 19 fill_sram_inverted $T=184 13148 1 0 $X=160 $Y=12432
XX73A2B172279_1 3 2 7 20 fill_sram_inverted $T=16 7916 1 0 $X=-8 $Y=7200
XX73A2B172279_2 3 2 7 20 fill_sram_inverted $T=184 7916 1 0 $X=160 $Y=7200
XX73A2B172281_1 3 2 8 21 fill_sram_inverted $T=16 10532 1 0 $X=-8 $Y=9816
XX73A2B172281_2 3 2 8 21 fill_sram_inverted $T=184 10532 1 0 $X=160 $Y=9816
XX73A2B172283_1 3 2 9 22 fill_sram_inverted $T=16 9224 1 0 $X=-8 $Y=8508
XX73A2B172283_2 3 2 9 22 fill_sram_inverted $T=184 9224 1 0 $X=160 $Y=8508
XX73A2B172285_1 3 2 10 23 fill_sram_inverted $T=16 1376 1 0 $X=-8 $Y=660
XX73A2B172285_2 3 2 10 23 fill_sram_inverted $T=184 1376 1 0 $X=160 $Y=660
XX73A2B172287_1 3 2 11 24 fill_sram_inverted $T=16 2684 1 0 $X=-8 $Y=1968
XX73A2B172287_2 3 2 11 24 fill_sram_inverted $T=184 2684 1 0 $X=160 $Y=1968
XX73A2B172289_1 3 2 12 25 fill_sram_inverted $T=16 3992 1 0 $X=-8 $Y=3276
XX73A2B172289_2 3 2 12 25 fill_sram_inverted $T=184 3992 1 0 $X=160 $Y=3276
XX73A2B172291_1 3 2 13 26 fill_sram_inverted $T=16 5300 1 0 $X=-8 $Y=4584
XX73A2B172291_2 3 2 13 26 fill_sram_inverted $T=184 5300 1 0 $X=160 $Y=4584
XX73A2B172293_1 3 2 14 27 fill_sram_inverted $T=16 6608 1 0 $X=-8 $Y=5892
XX73A2B172293_2 3 2 14 27 fill_sram_inverted $T=184 6608 1 0 $X=160 $Y=5892
XX73A2B172295_1 3 2 6 28 fill_sram $T=16 14458 0 0 $X=-8 $Y=14394
XX73A2B172295_2 3 2 6 28 fill_sram $T=184 14458 0 0 $X=160 $Y=14394
XX73A2B172297_1 3 2 5 19 fill_sram $T=16 11842 0 0 $X=-8 $Y=11778
XX73A2B172297_2 3 2 5 19 fill_sram $T=184 11842 0 0 $X=160 $Y=11778
XX73A2B172299_1 3 2 8 18 fill_sram $T=16 10534 0 0 $X=-8 $Y=10470
XX73A2B172299_2 3 2 8 18 fill_sram $T=184 10534 0 0 $X=160 $Y=10470
XX73A2B172301_1 3 2 14 20 fill_sram $T=16 6610 0 0 $X=-8 $Y=6546
XX73A2B172301_2 3 2 14 20 fill_sram $T=184 6610 0 0 $X=160 $Y=6546
XX73A2B172303_1 3 2 9 21 fill_sram $T=16 9226 0 0 $X=-8 $Y=9162
XX73A2B172303_2 3 2 9 21 fill_sram $T=184 9226 0 0 $X=160 $Y=9162
XX73A2B172305_1 3 2 7 22 fill_sram $T=16 7918 0 0 $X=-8 $Y=7854
XX73A2B172305_2 3 2 7 22 fill_sram $T=184 7918 0 0 $X=160 $Y=7854
XX73A2B172307_1 3 2 10 24 fill_sram $T=16 1378 0 0 $X=-8 $Y=1314
XX73A2B172307_2 3 2 10 24 fill_sram $T=184 1378 0 0 $X=160 $Y=1314
XX73A2B172309_1 3 2 11 25 fill_sram $T=16 2686 0 0 $X=-8 $Y=2622
XX73A2B172309_2 3 2 11 25 fill_sram $T=184 2686 0 0 $X=160 $Y=2622
XX73A2B172311_1 3 2 12 26 fill_sram $T=16 3994 0 0 $X=-8 $Y=3930
XX73A2B172311_2 3 2 12 26 fill_sram $T=184 3994 0 0 $X=160 $Y=3930
XX73A2B172313_1 3 2 13 27 fill_sram $T=16 5302 0 0 $X=-8 $Y=5238
XX73A2B172313_2 3 2 13 27 fill_sram $T=184 5302 0 0 $X=160 $Y=5238
XX73A2B172315_1 3 2 15 23 fill_sram $T=16 70 0 0 $X=-8 $Y=6
XX73A2B172315_2 3 2 15 23 fill_sram $T=184 70 0 0 $X=160 $Y=6
.ends sram_lvs_grid
.subckt sram_array_1r_4c 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22
XX73A2B172379 8 10 9 14 13 12 11 21 22 sram_6T_1finger $T=3024 16 0 0 $X=2970 $Y=-64
XX73A2B172380 6 10 7 16 15 12 11 21 22 sram_6T_1finger $T=2016 16 0 0 $X=1962 $Y=-64
XX73A2B172381 4 10 5 18 17 12 11 21 22 sram_6T_1finger $T=1008 16 0 0 $X=954 $Y=-64
XX73A2B172382 2 10 3 20 19 12 11 21 22 sram_6T_1finger $T=0 16 0 0 $X=-54 $Y=-64
XX73A2B172383 11 12 21 22 fill_sram $T=2826 0 0 0 $X=2802 $Y=-64
XX73A2B172384 11 12 21 22 fill_sram $T=1818 0 0 0 $X=1794 $Y=-64
XX73A2B172385 11 12 21 22 fill_sram $T=810 0 0 0 $X=786 $Y=-64
.ends sram_array_1r_4c
.subckt equalizer 2 3 4 5 6 7 8
XX73A2B172386_1 6 5 2 2 7 2 8 fill_sram_nmos $T=24 70 0 0 $X=0 $Y=6
XX73A2B172386_2 6 5 5 5 7 5 8 fill_sram_nmos $T=192 70 0 0 $X=168 $Y=6
XX73A2B172386_3 6 5 2 2 7 2 8 fill_sram_nmos $T=360 70 0 0 $X=335 $Y=6
XX73A2B172386_4 6 5 4 4 7 4 8 fill_sram_nmos $T=528 70 0 0 $X=504 $Y=6
XX73A2B172386_5 6 5 2 2 7 2 8 fill_sram_nmos $T=696 70 0 0 $X=672 $Y=6
XX73A2B172386_6 6 5 5 5 7 5 8 fill_sram_nmos $T=864 70 0 0 $X=840 $Y=6
XX73A2B172386_7 6 5 4 4 7 4 8 fill_sram_nmos $T=1032 70 0 0 $X=1008 $Y=6
XX73A2B172386_8 6 5 5 5 7 5 8 fill_sram_nmos $T=1200 70 0 0 $X=1176 $Y=6
.ends equalizer
.subckt buffer_top 2 3 4 5 6 7 8
XX73A2B172394 2 3 5 6 2 7 8 inverter_buf_top_level_v1 $T=504 86 0 0 $X=504 $Y=6
XX73A2B172395 4 3 5 6 7 8 inverter_buf_top_leve $T=0 86 0 0 $X=0 $Y=6
.ends buffer_top
.subckt column_decoder_read_cell 2 3 4 5 6 7 8 9 10 11 12
+	13
XX73A2B172396_1 9 8 12 2 13 fill_sram_inverted_pmos_read $T=24 716 1 0 $X=0 $Y=0
XX73A2B172396_2 9 8 12 10 13 fill_sram_inverted_pmos_read $T=192 716 1 0 $X=168 $Y=0
XX73A2B172396_3 9 8 12 7 13 fill_sram_inverted_pmos_read $T=360 716 1 0 $X=335 $Y=0
XX73A2B172396_4 9 8 12 11 13 fill_sram_inverted_pmos_read $T=528 716 1 0 $X=504 $Y=0
XX73A2B172396_5 9 8 12 5 13 fill_sram_inverted_pmos_read $T=696 716 1 0 $X=672 $Y=0
.ends column_decoder_read_cell
.subckt buffer_top_inverted 2 3 4 5 6 7 8
XX73A2B172401 2 3 5 6 2 7 8 inverter_buf_top_level_v1 $T=504 86 0 0 $X=504 $Y=6
XX73A2B172402 4 3 5 6 7 8 inverter_buf_top_leve $T=0 86 0 0 $X=0 $Y=6
.ends buffer_top_inverted
.subckt write_buffer_cell 4 6 7 8 11 12 13 14 15 18 19
MM1 8 3 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1848 $Y=864  $PIN_XY=1878,862,1848,864,1818,862 $DEVICE_ID=1001
MM2 3 9 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1848 $Y=390  $PIN_XY=1878,572,1848,390,1818,572 $DEVICE_ID=1001
MM3 11 6 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1680 $Y=390  $PIN_XY=1710,572,1680,390,1650,572 $DEVICE_ID=1001
MM4 16 4 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1512 $Y=390  $PIN_XY=1542,572,1512,390,1482,572 $DEVICE_ID=1001
MM5 11 4 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1176 $Y=390  $PIN_XY=1206,572,1176,390,1146,572 $DEVICE_ID=1001
MM6 10 5 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=840 $Y=390  $PIN_XY=870,572,840,390,810,572 $DEVICE_ID=1001
MM7 17 6 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=672 $Y=390  $PIN_XY=702,572,672,390,642,572 $DEVICE_ID=1001
MM8 11 2 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=504 $Y=864  $PIN_XY=534,862,504,864,474,862 $DEVICE_ID=1001
MM9 11 10 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=504 $Y=390  $PIN_XY=534,572,504,390,474,572 $DEVICE_ID=1001
XX73A2B172403 4 5 11 12 14 15 18 inverter_write $T=1398 700 0 180 $X=954 $Y=0
XX73A2B172404_1 11 13 14 19 fill_sram $T=642 718 0 0 $X=618 $Y=653
XX73A2B172404_2 11 13 14 19 fill_sram $T=810 718 0 0 $X=786 $Y=653
XX73A2B172404_3 11 13 14 19 fill_sram $T=978 718 0 0 $X=954 $Y=653
XX73A2B172404_4 11 13 14 19 fill_sram $T=1146 718 0 0 $X=1122 $Y=653
XX73A2B172404_5 11 13 14 19 fill_sram $T=1314 718 0 0 $X=1290 $Y=653
XX73A2B172404_6 11 13 14 19 fill_sram $T=1482 718 0 0 $X=1458 $Y=653
XX73A2B172410_1 13 11 14 8 19 fill_sram_inverted_pmos_write $T=2046 718 1 180 $X=1794 $Y=653
XX73A2B172410_2 13 11 14 11 19 fill_sram_inverted_pmos_write $T=1878 718 1 180 $X=1626 $Y=653
XX73A2B172412_1 13 11 14 7 19 fill_sram_inverted_pmos_write $T=306 718 0 0 $X=282 $Y=653
XX73A2B172412_2 13 11 14 11 19 fill_sram_inverted_pmos_write $T=474 718 0 0 $X=450 $Y=653
XX73A2B172414 9 3 4 6 12 11 16 14 15 18 and_v1 $T=1344 716 1 0 $X=1290 $Y=0
XX73A2B172415 10 2 5 6 12 11 17 14 15 18 and $T=1008 716 0 180 $X=282 $Y=0
.ends write_buffer_cell
.subckt column_decoder_write_cell 2 3 4 5 6 7 8 9 10
XX73A2B172416_1 8 7 9 10 fill_sram_inverted_write_pmos $T=24 70 0 0 $X=0 $Y=6
XX73A2B172416_2 8 7 9 10 fill_sram_inverted_write_pmos $T=192 70 0 0 $X=168 $Y=6
XX73A2B172416_3 8 7 9 10 fill_sram_inverted_write_pmos $T=360 70 0 0 $X=335 $Y=6
XX73A2B172416_4 8 7 9 10 fill_sram_inverted_write_pmos $T=528 70 0 0 $X=504 $Y=6
.ends column_decoder_write_cell
.subckt VCELLR3 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 23
MM1 3 13 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1230 $Y=1524  $PIN_XY=1260,1522,1230,1524,1200,1522 $DEVICE_ID=1001
MM2 3 11 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=1524  $PIN_XY=924,1522,894,1524,864,1522 $DEVICE_ID=1001
MM3 3 9 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=558 $Y=1524  $PIN_XY=588,1522,558,1524,528,1522 $DEVICE_ID=1001
MM4 3 6 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=1524  $PIN_XY=252,1522,222,1524,192,1522 $DEVICE_ID=1001
MM5 3 7 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=222 $Y=2232  $PIN_XY=(252,2346,252,2176),222,2232,(192,2346,192,2176) $DEVICE_ID=1003
MM6 2 5 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=222 $Y=924  $PIN_XY=(252,1038,252,868),222,924,(192,1038,192,868) $DEVICE_ID=1003
XX73A2B172420_1 16 15 19 22 fill_sram_inverted $T=360 1376 1 0 $X=335 $Y=660
XX73A2B172420_2 16 15 19 22 fill_sram_inverted $T=528 1376 1 0 $X=504 $Y=660
XX73A2B172420_3 16 15 19 22 fill_sram_inverted $T=696 1376 1 0 $X=672 $Y=660
XX73A2B172420_4 16 15 19 22 fill_sram_inverted $T=864 1376 1 0 $X=840 $Y=660
XX73A2B172420_5 16 15 19 22 fill_sram_inverted $T=1032 1376 1 0 $X=1008 $Y=660
XX73A2B172420_6 16 15 19 22 fill_sram_inverted $T=1200 1376 1 0 $X=1176 $Y=660
XX73A2B172426_1 18 17 20 23 fill_sram_inverted $T=360 2684 1 0 $X=335 $Y=1968
XX73A2B172426_2 18 17 20 23 fill_sram_inverted $T=528 2684 1 0 $X=504 $Y=1968
XX73A2B172426_3 18 17 20 23 fill_sram_inverted $T=696 2684 1 0 $X=672 $Y=1968
XX73A2B172426_4 18 17 20 23 fill_sram_inverted $T=864 2684 1 0 $X=840 $Y=1968
XX73A2B172426_5 18 17 20 23 fill_sram_inverted $T=1032 2684 1 0 $X=1008 $Y=1968
XX73A2B172426_6 18 17 20 23 fill_sram_inverted $T=1200 2684 1 0 $X=1176 $Y=1968
XX73A2B172432_1 16 15 19 22 fill_sram_inverted_nmos $T=24 1376 1 0 $X=24 $Y=660
XX73A2B172432_2 16 15 19 22 fill_sram_inverted_nmos $T=192 1376 1 0 $X=192 $Y=660
XX73A2B172434_1 18 17 20 23 fill_sram_inverted_nmos $T=24 2684 1 0 $X=24 $Y=1968
XX73A2B172434_2 18 17 20 23 fill_sram_inverted_nmos $T=192 2684 1 0 $X=192 $Y=1968
XX73A2B172436_1 15 14 21 14 22 fill_sram_pmos $T=24 70 0 0 $X=24 $Y=6
XX73A2B172436_2 15 14 21 2 22 fill_sram_pmos $T=192 70 0 0 $X=192 $Y=6
XX73A2B172436_3 15 14 21 14 22 fill_sram_pmos $T=360 70 0 0 $X=360 $Y=6
XX73A2B172436_4 15 14 21 2 22 fill_sram_pmos $T=528 70 0 0 $X=528 $Y=6
XX73A2B172436_5 15 14 21 14 22 fill_sram_pmos $T=696 70 0 0 $X=696 $Y=6
XX73A2B172436_6 15 14 21 2 22 fill_sram_pmos $T=864 70 0 0 $X=864 $Y=6
XX73A2B172436_7 15 14 21 14 22 fill_sram_pmos $T=1032 70 0 0 $X=1032 $Y=6
XX73A2B172436_8 15 14 21 2 22 fill_sram_pmos $T=1200 70 0 0 $X=1200 $Y=6
XX73A2B172444_1 17 16 19 16 23 fill_sram_pmos $T=24 1378 0 0 $X=24 $Y=1314
XX73A2B172444_2 17 16 19 3 23 fill_sram_pmos $T=192 1378 0 0 $X=192 $Y=1314
XX73A2B172444_3 17 16 19 16 23 fill_sram_pmos $T=360 1378 0 0 $X=360 $Y=1314
XX73A2B172444_4 17 16 19 3 23 fill_sram_pmos $T=528 1378 0 0 $X=528 $Y=1314
XX73A2B172444_5 17 16 19 16 23 fill_sram_pmos $T=696 1378 0 0 $X=696 $Y=1314
XX73A2B172444_6 17 16 19 3 23 fill_sram_pmos $T=864 1378 0 0 $X=864 $Y=1314
XX73A2B172444_7 17 16 19 16 23 fill_sram_pmos $T=1032 1378 0 0 $X=1032 $Y=1314
XX73A2B172444_8 17 16 19 3 23 fill_sram_pmos $T=1200 1378 0 0 $X=1200 $Y=1314
.ends VCELLR3

* Hierarchy Level 2
.subckt bitline_conditioning 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 23
+	24
MM1 18 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=7728 $Y=419  $PIN_XY=(7758,508,7758,338),7728,419,(7698,508,7698,338) $DEVICE_ID=1003
MM2 20 2 18 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=7560 $Y=419  $PIN_XY=(7590,508,7590,338),7560,419,(7530,508,7530,338) $DEVICE_ID=1003
MM3 18 2 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=7392 $Y=419  $PIN_XY=(7422,508,7422,338),7392,419,(7362,508,7362,338) $DEVICE_ID=1003
MM4 16 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=7224 $Y=887  $PIN_XY=(7254,968,7254,798),7224,887,(7194,968,7194,798) $DEVICE_ID=1003
MM5 17 2 18 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=7224 $Y=419  $PIN_XY=(7254,508,7254,338),7224,419,(7194,508,7194,338) $DEVICE_ID=1003
MM6 20 2 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=7056 $Y=887  $PIN_XY=(7086,968,7086,798),7056,887,(7026,968,7026,798) $DEVICE_ID=1003
MM7 16 2 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=6888 $Y=887  $PIN_XY=(6918,968,6918,798),6888,887,(6858,968,6858,798) $DEVICE_ID=1003
MM8 20 2 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=6888 $Y=419  $PIN_XY=(6918,508,6918,338),6888,419,(6858,508,6858,338) $DEVICE_ID=1003
MM9 15 2 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=6720 $Y=887  $PIN_XY=(6750,968,6750,798),6720,887,(6690,968,6690,798) $DEVICE_ID=1003
MM10 17 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=6720 $Y=419  $PIN_XY=(6750,508,6750,338),6720,419,(6690,508,6690,338) $DEVICE_ID=1003
MM11 20 2 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=6384 $Y=887  $PIN_XY=(6414,968,6414,798),6384,887,(6354,968,6354,798) $DEVICE_ID=1003
MM12 15 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=6216 $Y=887  $PIN_XY=(6246,968,6246,798),6216,887,(6186,968,6186,798) $DEVICE_ID=1003
MM13 14 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=5712 $Y=419  $PIN_XY=(5742,508,5742,338),5712,419,(5682,508,5682,338) $DEVICE_ID=1003
MM14 20 2 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=5544 $Y=419  $PIN_XY=(5574,508,5574,338),5544,419,(5514,508,5514,338) $DEVICE_ID=1003
MM15 14 2 13 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=5376 $Y=419  $PIN_XY=(5406,508,5406,338),5376,419,(5346,508,5346,338) $DEVICE_ID=1003
MM16 12 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=5208 $Y=887  $PIN_XY=(5238,968,5238,798),5208,887,(5178,968,5178,798) $DEVICE_ID=1003
MM17 13 2 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=5208 $Y=419  $PIN_XY=(5238,508,5238,338),5208,419,(5178,508,5178,338) $DEVICE_ID=1003
MM18 20 2 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=5040 $Y=887  $PIN_XY=(5070,968,5070,798),5040,887,(5010,968,5010,798) $DEVICE_ID=1003
MM19 12 2 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=4872 $Y=887  $PIN_XY=(4902,968,4902,798),4872,887,(4842,968,4842,798) $DEVICE_ID=1003
MM20 20 2 13 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=4872 $Y=419  $PIN_XY=(4902,508,4902,338),4872,419,(4842,508,4842,338) $DEVICE_ID=1003
MM21 11 2 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=4704 $Y=887  $PIN_XY=(4734,968,4734,798),4704,887,(4674,968,4674,798) $DEVICE_ID=1003
MM22 13 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=4704 $Y=419  $PIN_XY=(4734,508,4734,338),4704,419,(4674,508,4674,338) $DEVICE_ID=1003
MM23 20 2 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=4368 $Y=887  $PIN_XY=(4398,968,4398,798),4368,887,(4338,968,4338,798) $DEVICE_ID=1003
MM24 11 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=4200 $Y=887  $PIN_XY=(4230,968,4230,798),4200,887,(4170,968,4170,798) $DEVICE_ID=1003
MM25 10 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3696 $Y=419  $PIN_XY=(3726,508,3726,338),3696,419,(3666,508,3666,338) $DEVICE_ID=1003
MM26 20 2 10 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3528 $Y=419  $PIN_XY=(3558,508,3558,338),3528,419,(3498,508,3498,338) $DEVICE_ID=1003
MM27 10 2 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3360 $Y=419  $PIN_XY=(3390,508,3390,338),3360,419,(3330,508,3330,338) $DEVICE_ID=1003
MM28 8 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3192 $Y=887  $PIN_XY=(3222,968,3222,798),3192,887,(3162,968,3162,798) $DEVICE_ID=1003
MM29 9 2 10 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=419  $PIN_XY=(3222,508,3222,338),3192,419,(3162,508,3162,338) $DEVICE_ID=1003
MM30 20 2 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3024 $Y=887  $PIN_XY=(3054,968,3054,798),3024,887,(2994,968,2994,798) $DEVICE_ID=1003
MM31 8 2 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=2856 $Y=887  $PIN_XY=(2886,968,2886,798),2856,887,(2826,968,2826,798) $DEVICE_ID=1003
MM32 20 2 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=2856 $Y=419  $PIN_XY=(2886,508,2886,338),2856,419,(2826,508,2826,338) $DEVICE_ID=1003
MM33 7 2 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=2688 $Y=887  $PIN_XY=(2718,968,2718,798),2688,887,(2658,968,2658,798) $DEVICE_ID=1003
MM34 9 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=2688 $Y=419  $PIN_XY=(2718,508,2718,338),2688,419,(2658,508,2658,338) $DEVICE_ID=1003
MM35 20 2 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=2352 $Y=887  $PIN_XY=(2382,968,2382,798),2352,887,(2322,968,2322,798) $DEVICE_ID=1003
MM36 7 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=2184 $Y=887  $PIN_XY=(2214,968,2214,798),2184,887,(2154,968,2154,798) $DEVICE_ID=1003
MM37 6 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=1680 $Y=419  $PIN_XY=(1710,508,1710,338),1680,419,(1650,508,1650,338) $DEVICE_ID=1003
MM38 20 2 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=1512 $Y=419  $PIN_XY=(1542,508,1542,338),1512,419,(1482,508,1482,338) $DEVICE_ID=1003
MM39 6 2 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=1344 $Y=419  $PIN_XY=(1374,508,1374,338),1344,419,(1314,508,1314,338) $DEVICE_ID=1003
MM40 4 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=1176 $Y=887  $PIN_XY=(1206,968,1206,798),1176,887,(1146,968,1146,798) $DEVICE_ID=1003
MM41 5 2 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=1176 $Y=419  $PIN_XY=(1206,508,1206,338),1176,419,(1146,508,1146,338) $DEVICE_ID=1003
MM42 20 2 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=1008 $Y=887  $PIN_XY=(1038,968,1038,798),1008,887,(978,968,978,798) $DEVICE_ID=1003
MM43 4 2 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=840 $Y=887  $PIN_XY=(870,968,870,798),840,887,(810,968,810,798) $DEVICE_ID=1003
MM44 20 2 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=840 $Y=419  $PIN_XY=(870,508,870,338),840,419,(810,508,810,338) $DEVICE_ID=1003
MM45 3 2 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=672 $Y=887  $PIN_XY=(702,968,702,798),672,887,(642,968,642,798) $DEVICE_ID=1003
MM46 5 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=672 $Y=419  $PIN_XY=(702,508,702,338),672,419,(642,508,642,338) $DEVICE_ID=1003
MM47 20 2 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=336 $Y=887  $PIN_XY=(366,968,366,798),336,887,(306,968,306,798) $DEVICE_ID=1003
MM48 3 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=168 $Y=887  $PIN_XY=(198,968,198,798),168,887,(138,968,138,798) $DEVICE_ID=1003
XX73A2B172179_1 19 20 22 24 fill_sram $T=5850 0 0 0 $X=5826 $Y=-64
XX73A2B172179_2 19 20 22 24 fill_sram $T=6018 0 0 0 $X=5994 $Y=-64
XX73A2B172179_3 19 20 22 24 fill_sram $T=6186 0 0 0 $X=6162 $Y=-64
XX73A2B172179_4 19 20 22 24 fill_sram $T=6354 0 0 0 $X=6330 $Y=-64
XX73A2B172183_1 19 20 22 24 fill_sram $T=1818 0 0 0 $X=1794 $Y=-64
XX73A2B172183_2 19 20 22 24 fill_sram $T=1986 0 0 0 $X=1962 $Y=-64
XX73A2B172183_3 19 20 22 24 fill_sram $T=2154 0 0 0 $X=2130 $Y=-64
XX73A2B172183_4 19 20 22 24 fill_sram $T=2322 0 0 0 $X=2298 $Y=-64
XX73A2B172187_1 19 20 22 24 fill_sram $T=-30 0 0 0 $X=-54 $Y=-64
XX73A2B172187_2 19 20 22 24 fill_sram $T=138 0 0 0 $X=114 $Y=-64
XX73A2B172187_3 19 20 22 24 fill_sram $T=306 0 0 0 $X=282 $Y=-64
XX73A2B172190_1 19 20 22 24 fill_sram $T=3834 0 0 0 $X=3810 $Y=-64
XX73A2B172190_2 19 20 22 24 fill_sram $T=4002 0 0 0 $X=3977 $Y=-64
XX73A2B172190_3 19 20 22 24 fill_sram $T=4170 0 0 0 $X=4146 $Y=-64
XX73A2B172190_4 19 20 22 24 fill_sram $T=4338 0 0 0 $X=4314 $Y=-64
XX73A2B172194 14 2 13 20 19 22 24 equalizer $T=5934 -70 1 180 $X=4482 $Y=-64
XX73A2B172195 16 2 15 20 21 23 24 equalizer $T=7446 1376 0 180 $X=5994 $Y=590
XX73A2B172196 10 2 9 20 19 22 24 equalizer $T=3918 -70 1 180 $X=2466 $Y=-64
XX73A2B172197 8 2 7 20 21 23 24 equalizer $T=3414 1376 0 180 $X=1962 $Y=590
XX73A2B172198 12 2 11 20 21 23 24 equalizer $T=5430 1376 0 180 $X=3977 $Y=590
XX73A2B172199 6 2 5 20 19 22 24 equalizer $T=1902 -70 1 180 $X=450 $Y=-64
XX73A2B172200 4 2 3 20 21 23 24 equalizer $T=1398 1376 0 180 $X=-53 $Y=590
XX73A2B172201 18 2 17 20 19 22 24 equalizer $T=7950 -70 1 180 $X=6498 $Y=-64
XX73A2B172202_1 21 20 23 24 fill_sram_inverted $T=3330 1306 1 0 $X=3306 $Y=590
XX73A2B172202_2 21 20 23 24 fill_sram_inverted $T=3498 1306 1 0 $X=3474 $Y=590
XX73A2B172202_3 21 20 23 24 fill_sram_inverted $T=3666 1306 1 0 $X=3642 $Y=590
XX73A2B172202_4 21 20 23 24 fill_sram_inverted $T=3834 1306 1 0 $X=3810 $Y=590
XX73A2B172206_1 21 20 23 24 fill_sram_inverted $T=1314 1306 1 0 $X=1290 $Y=590
XX73A2B172206_2 21 20 23 24 fill_sram_inverted $T=1482 1306 1 0 $X=1458 $Y=590
XX73A2B172206_3 21 20 23 24 fill_sram_inverted $T=1650 1306 1 0 $X=1626 $Y=590
XX73A2B172206_4 21 20 23 24 fill_sram_inverted $T=1818 1306 1 0 $X=1794 $Y=590
XX73A2B172210_1 21 20 23 24 fill_sram_inverted $T=7362 1306 1 0 $X=7338 $Y=590
XX73A2B172210_2 21 20 23 24 fill_sram_inverted $T=7530 1306 1 0 $X=7506 $Y=590
XX73A2B172210_3 21 20 23 24 fill_sram_inverted $T=7698 1306 1 0 $X=7674 $Y=590
XX73A2B172213_1 21 20 23 24 fill_sram_inverted $T=5346 1306 1 0 $X=5322 $Y=590
XX73A2B172213_2 21 20 23 24 fill_sram_inverted $T=5514 1306 1 0 $X=5490 $Y=590
XX73A2B172213_3 21 20 23 24 fill_sram_inverted $T=5682 1306 1 0 $X=5658 $Y=590
XX73A2B172213_4 21 20 23 24 fill_sram_inverted $T=5850 1306 1 0 $X=5826 $Y=590
.ends bitline_conditioning
.subckt buffer_array 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17
MM1 10 2 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6774 $Y=396  $PIN_XY=6804,214,6774,396,6744,214 $DEVICE_ID=1001
MM2 12 2 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6606 $Y=396  $PIN_XY=6636,214,6606,396,6576,214 $DEVICE_ID=1001
MM3 10 3 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6270 $Y=396  $PIN_XY=6300,214,6270,396,6240,214 $DEVICE_ID=1001
MM4 2 3 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6102 $Y=396  $PIN_XY=6132,214,6102,396,6072,214 $DEVICE_ID=1001
MM5 10 4 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4758 $Y=396  $PIN_XY=4788,214,4758,396,4728,214 $DEVICE_ID=1001
MM6 13 4 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4590 $Y=396  $PIN_XY=4620,214,4590,396,4560,214 $DEVICE_ID=1001
MM7 10 5 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4254 $Y=396  $PIN_XY=4284,214,4254,396,4224,214 $DEVICE_ID=1001
MM8 4 5 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4086 $Y=396  $PIN_XY=4116,214,4086,396,4056,214 $DEVICE_ID=1001
MM9 10 6 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2742 $Y=396  $PIN_XY=2772,214,2742,396,2712,214 $DEVICE_ID=1001
MM10 14 6 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2574 $Y=396  $PIN_XY=2604,214,2574,396,2544,214 $DEVICE_ID=1001
MM11 10 7 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2238 $Y=396  $PIN_XY=2268,214,2238,396,2208,214 $DEVICE_ID=1001
MM12 6 7 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2070 $Y=396  $PIN_XY=2100,214,2070,396,2040,214 $DEVICE_ID=1001
MM13 10 8 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=894 $Y=396  $PIN_XY=924,214,894,396,864,214 $DEVICE_ID=1001
MM14 15 8 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=726 $Y=396  $PIN_XY=756,214,726,396,696,214 $DEVICE_ID=1001
MM15 10 9 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=396  $PIN_XY=420,214,390,396,360,214 $DEVICE_ID=1001
MM16 8 9 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=396  $PIN_XY=252,214,222,396,192,214 $DEVICE_ID=1001
XX73A2B172217 12 2 3 10 11 16 17 buffer_top $T=5880 0 0 0 $X=5880 $Y=6
XX73A2B172218 13 4 5 10 11 16 17 buffer_top $T=3864 0 0 0 $X=3864 $Y=6
XX73A2B172219 14 6 7 10 11 16 17 buffer_top $T=1848 0 0 0 $X=1848 $Y=6
XX73A2B172220 15 8 9 10 11 16 17 buffer_top $T=0 0 0 0 $X=0 $Y=6
XX73A2B172221_1 10 11 16 17 fill_sram $T=6912 70 0 0 $X=6888 $Y=6
XX73A2B172221_2 10 11 16 17 fill_sram $T=7080 70 0 0 $X=7056 $Y=6
XX73A2B172223_1 10 11 16 17 fill_sram $T=4896 70 0 0 $X=4872 $Y=6
XX73A2B172223_2 10 11 16 17 fill_sram $T=5064 70 0 0 $X=5040 $Y=6
XX73A2B172223_3 10 11 16 17 fill_sram $T=5232 70 0 0 $X=5208 $Y=6
XX73A2B172223_4 10 11 16 17 fill_sram $T=5400 70 0 0 $X=5376 $Y=6
XX73A2B172223_5 10 11 16 17 fill_sram $T=5568 70 0 0 $X=5544 $Y=6
XX73A2B172223_6 10 11 16 17 fill_sram $T=5736 70 0 0 $X=5712 $Y=6
XX73A2B172229_1 10 11 16 17 fill_sram $T=1032 70 0 0 $X=1008 $Y=6
XX73A2B172229_2 10 11 16 17 fill_sram $T=1200 70 0 0 $X=1176 $Y=6
XX73A2B172229_3 10 11 16 17 fill_sram $T=1368 70 0 0 $X=1344 $Y=6
XX73A2B172229_4 10 11 16 17 fill_sram $T=1536 70 0 0 $X=1512 $Y=6
XX73A2B172229_5 10 11 16 17 fill_sram $T=1704 70 0 0 $X=1680 $Y=6
XX73A2B172234_1 10 11 16 17 fill_sram $T=2880 70 0 0 $X=2856 $Y=6
XX73A2B172234_2 10 11 16 17 fill_sram $T=3048 70 0 0 $X=3024 $Y=6
XX73A2B172234_3 10 11 16 17 fill_sram $T=3216 70 0 0 $X=3192 $Y=6
XX73A2B172234_4 10 11 16 17 fill_sram $T=3384 70 0 0 $X=3360 $Y=6
XX73A2B172234_5 10 11 16 17 fill_sram $T=3552 70 0 0 $X=3528 $Y=6
XX73A2B172234_6 10 11 16 17 fill_sram $T=3720 70 0 0 $X=3696 $Y=6
.ends buffer_array
.subckt column_decoder_read 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 23
+	24 25 26 27 28
XX73A2B172240 4 2 3 5 6 7 18 17 21 22 19 
+	20 column_decoder_read_cell $T=7564 0 0 0 $X=7564 $Y=0
XX73A2B172241 8 2 3 9 6 10 18 17 23 24 19 
+	20 column_decoder_read_cell $T=5548 0 0 0 $X=5548 $Y=0
XX73A2B172242 11 2 3 12 6 13 18 17 25 26 19 
+	20 column_decoder_read_cell $T=3532 0 0 0 $X=3532 $Y=0
XX73A2B172243 14 2 3 15 6 16 18 17 27 28 19 
+	20 column_decoder_read_cell $T=1684 0 0 0 $X=1684 $Y=0
XX73A2B172244_1 18 17 19 20 fill_sram_inverted_read $T=8428 716 1 0 $X=8404 $Y=0
XX73A2B172244_2 18 17 19 20 fill_sram_inverted_read $T=8596 716 1 0 $X=8572 $Y=0
XX73A2B172244_3 18 17 19 20 fill_sram_inverted_read $T=8764 716 1 0 $X=8740 $Y=0
XX73A2B172247_1 18 17 19 20 fill_sram_inverted_read $T=6412 716 1 0 $X=6388 $Y=0
XX73A2B172247_2 18 17 19 20 fill_sram_inverted_read $T=6580 716 1 0 $X=6556 $Y=0
XX73A2B172247_3 18 17 19 20 fill_sram_inverted_read $T=6748 716 1 0 $X=6724 $Y=0
XX73A2B172247_4 18 17 19 20 fill_sram_inverted_read $T=6916 716 1 0 $X=6892 $Y=0
XX73A2B172247_5 18 17 19 20 fill_sram_inverted_read $T=7084 716 1 0 $X=7060 $Y=0
XX73A2B172247_6 18 17 19 20 fill_sram_inverted_read $T=7252 716 1 0 $X=7228 $Y=0
XX73A2B172247_7 18 17 19 20 fill_sram_inverted_read $T=7420 716 1 0 $X=7396 $Y=0
XX73A2B172254_1 18 17 19 20 fill_sram_inverted_read $T=4396 716 1 0 $X=4372 $Y=0
XX73A2B172254_2 18 17 19 20 fill_sram_inverted_read $T=4564 716 1 0 $X=4540 $Y=0
XX73A2B172254_3 18 17 19 20 fill_sram_inverted_read $T=4732 716 1 0 $X=4708 $Y=0
XX73A2B172254_4 18 17 19 20 fill_sram_inverted_read $T=4900 716 1 0 $X=4876 $Y=0
XX73A2B172254_5 18 17 19 20 fill_sram_inverted_read $T=5068 716 1 0 $X=5044 $Y=0
XX73A2B172254_6 18 17 19 20 fill_sram_inverted_read $T=5236 716 1 0 $X=5212 $Y=0
XX73A2B172254_7 18 17 19 20 fill_sram_inverted_read $T=5404 716 1 0 $X=5380 $Y=0
XX73A2B172261_1 18 17 19 20 fill_sram_inverted_read $T=2548 716 1 0 $X=2524 $Y=0
XX73A2B172261_2 18 17 19 20 fill_sram_inverted_read $T=2716 716 1 0 $X=2692 $Y=0
XX73A2B172261_3 18 17 19 20 fill_sram_inverted_read $T=2884 716 1 0 $X=2860 $Y=0
XX73A2B172261_4 18 17 19 20 fill_sram_inverted_read $T=3052 716 1 0 $X=3028 $Y=0
XX73A2B172261_5 18 17 19 20 fill_sram_inverted_read $T=3220 716 1 0 $X=3196 $Y=0
XX73A2B172261_6 18 17 19 20 fill_sram_inverted_read $T=3388 716 1 0 $X=3364 $Y=0
XX73A2B172267_1 18 17 19 20 fill_sram_inverted_read $T=1036 716 1 0 $X=1012 $Y=0
XX73A2B172267_2 18 17 19 20 fill_sram_inverted_read $T=1204 716 1 0 $X=1180 $Y=0
XX73A2B172267_3 18 17 19 20 fill_sram_inverted_read $T=1372 716 1 0 $X=1348 $Y=0
XX73A2B172267_4 18 17 19 20 fill_sram_inverted_read $T=1540 716 1 0 $X=1516 $Y=0
.ends column_decoder_read
.subckt row_decoder_4_16 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 23
+	24 25 26 27 28 29 30 31 32 33 34
+	35 36 37 38 39 40 41 42 43 44 45
+	46 47 48 49 50 51 52 53 54 55 56
+	57 58 59 60 61 62
MM1 43 6 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2520 $Y=10790  $PIN_XY=2550,10608,2520,10790,2490,10608 $DEVICE_ID=1001
MM2 25 10 36 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2520 $Y=7994  $PIN_XY=2550,7992,2520,7994,2490,7992 $DEVICE_ID=1001
MM3 21 10 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2520 $Y=5378  $PIN_XY=2550,5376,2520,5378,2490,5376 $DEVICE_ID=1001
MM4 16 6 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2520 $Y=2762  $PIN_XY=2550,2760,2520,2762,2490,2760 $DEVICE_ID=1001
MM5 10 6 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2352 $Y=10790  $PIN_XY=2382,10608,2352,10790,2322,10608 $DEVICE_ID=1001
MM6 25 9 36 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2184 $Y=7994  $PIN_XY=2214,7992,2184,7994,2154,7992 $DEVICE_ID=1001
MM7 21 5 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2184 $Y=5378  $PIN_XY=2214,5376,2184,5378,2154,5376 $DEVICE_ID=1001
MM8 16 9 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2184 $Y=2762  $PIN_XY=2214,2760,2184,2762,2154,2760 $DEVICE_ID=1001
MM9 43 5 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1848 $Y=10790  $PIN_XY=1878,10608,1848,10790,1818,10608 $DEVICE_ID=1001
MM10 25 3 36 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1848 $Y=7994  $PIN_XY=1878,7992,1848,7994,1818,7992 $DEVICE_ID=1001
MM11 21 3 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1848 $Y=5378  $PIN_XY=1878,5376,1848,5378,1818,5376 $DEVICE_ID=1001
MM12 16 3 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1848 $Y=2762  $PIN_XY=1878,2760,1848,2762,1818,2760 $DEVICE_ID=1001
MM13 9 5 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1680 $Y=10790  $PIN_XY=1710,10608,1680,10790,1650,10608 $DEVICE_ID=1001
MM14 25 4 36 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1512 $Y=7994  $PIN_XY=1542,7992,1512,7994,1482,7992 $DEVICE_ID=1001
MM15 21 4 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1512 $Y=5378  $PIN_XY=1542,5376,1512,5378,1482,5376 $DEVICE_ID=1001
MM16 16 4 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1512 $Y=2762  $PIN_XY=1542,2760,1512,2762,1482,2760 $DEVICE_ID=1001
MM17 23 10 36 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1176 $Y=7994  $PIN_XY=1206,7992,1176,7994,1146,7992 $DEVICE_ID=1001
MM18 18 10 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1176 $Y=5378  $PIN_XY=1206,5376,1176,5378,1146,5376 $DEVICE_ID=1001
MM19 13 6 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1176 $Y=2762  $PIN_XY=1206,2760,1176,2762,1146,2760 $DEVICE_ID=1001
MM20 43 3 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1008 $Y=10790  $PIN_XY=1038,10608,1008,10790,978,10608 $DEVICE_ID=1001
MM21 8 3 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=840 $Y=10790  $PIN_XY=870,10608,840,10790,810,10608 $DEVICE_ID=1001
MM22 23 9 36 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=840 $Y=7994  $PIN_XY=870,7992,840,7994,810,7992 $DEVICE_ID=1001
MM23 18 5 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=840 $Y=5378  $PIN_XY=870,5376,840,5378,810,5376 $DEVICE_ID=1001
MM24 13 9 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=840 $Y=2762  $PIN_XY=870,2760,840,2762,810,2760 $DEVICE_ID=1001
MM25 23 3 36 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=504 $Y=7994  $PIN_XY=534,7992,504,7994,474,7992 $DEVICE_ID=1001
MM26 18 3 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=504 $Y=5378  $PIN_XY=534,5376,504,5378,474,5376 $DEVICE_ID=1001
MM27 13 3 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=504 $Y=2762  $PIN_XY=534,2760,504,2762,474,2760 $DEVICE_ID=1001
MM28 43 4 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=336 $Y=10790  $PIN_XY=366,10608,336,10790,306,10608 $DEVICE_ID=1001
MM29 7 4 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=10790  $PIN_XY=198,10608,168,10790,138,10608 $DEVICE_ID=1001
MM30 23 7 36 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=168 $Y=7994  $PIN_XY=198,7992,168,7994,138,7992 $DEVICE_ID=1001
MM31 18 7 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=168 $Y=5378  $PIN_XY=198,5376,168,5378,138,5376 $DEVICE_ID=1001
MM32 13 7 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=168 $Y=2762  $PIN_XY=198,2760,168,2762,138,2760 $DEVICE_ID=1001
XX73A2B172317 11 12 7 2 7 2 3 8 5 5 6 
+	6 28 29 30 31 27 45 46 47 54 55 VCELLR3 $T=-54 -70 0 0 $X=-54 $Y=-64
XX73A2B172318 13 17 7 2 7 2 3 8 9 9 6 
+	6 27 33 34 35 32 48 49 46 56 57 VCELLR3 $T=-54 2546 0 0 $X=-54 $Y=2552
XX73A2B172319 18 19 7 2 7 2 3 8 5 5 10 
+	10 32 37 38 39 36 50 51 49 58 59 VCELLR3 $T=-54 5162 0 0 $X=-54 $Y=5168
XX73A2B172320 23 24 7 2 7 2 3 8 9 9 10 
+	10 36 40 41 42 43 52 53 51 60 61 VCELLR3 $T=-54 7778 0 0 $X=-54 $Y=7784
XX73A2B172321 14 15 4 2 4 2 3 8 5 5 6 
+	6 28 29 30 31 27 45 46 47 54 55 VCELLR3 $T=1290 -70 0 0 $X=1290 $Y=-64
XX73A2B172322 16 20 4 2 4 2 3 8 9 9 6 
+	6 27 33 34 35 32 48 49 46 56 57 VCELLR3 $T=1290 2546 0 0 $X=1290 $Y=2552
XX73A2B172323 21 22 4 2 4 2 3 8 5 5 10 
+	10 32 37 38 39 36 50 51 49 58 59 VCELLR3 $T=1290 5162 0 0 $X=1290 $Y=5168
XX73A2B172324 25 26 4 2 4 2 3 8 9 9 10 
+	10 36 40 41 42 43 52 53 51 60 61 VCELLR3 $T=1290 7778 0 0 $X=1290 $Y=7784
XX73A2B172325 43 44 53 62 fill_sram $T=474 10464 0 0 $X=450 $Y=10400
XX73A2B172326 43 44 53 62 fill_sram $T=1986 10464 0 0 $X=1962 $Y=10400
XX73A2B172327_1 43 44 53 62 fill_sram $T=1146 10464 0 0 $X=1122 $Y=10400
XX73A2B172327_2 43 44 53 62 fill_sram $T=1314 10464 0 0 $X=1290 $Y=10400
XX73A2B172329 8 3 43 44 53 62 inverter_row_decoder $T=618 10480 0 0 $X=618 $Y=10400
XX73A2B172330 10 6 43 44 53 62 inverter_row_decoder $T=2130 10480 0 0 $X=2130 $Y=10400
XX73A2B172331 9 5 43 44 53 62 inverter_row_decoder $T=1458 10480 0 0 $X=1458 $Y=10400
XX73A2B172332 7 4 43 44 53 62 inverter_row_decoder $T=-54 10480 0 0 $X=-54 $Y=10400
.ends row_decoder_4_16
.subckt column_decoder_write 2 4 5 6 7 8 9 10 11 12 13
+	14 15 16 17 18 19 20 21 22 23 24
+	25 26 27 28 29 30 31 32 33 34 35
+	36 37 38 39 40 41 42
MM1 34 13 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=336 $Y=1704  $PIN_XY=366,1522,336,1704,306,1522 $DEVICE_ID=1001
MM2 34 2 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=336 $Y=1050  $PIN_XY=366,1232,336,1050,306,1232 $DEVICE_ID=1001
MM3 3 13 34 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=1704  $PIN_XY=198,1522,168,1704,138,1522 $DEVICE_ID=1001
MM4 4 2 34 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=1050  $PIN_XY=198,1232,168,1050,138,1232 $DEVICE_ID=1001
MM5 35 13 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=336 $Y=1704  $PIN_XY=(366,1886,366,1716),336,1704,(306,1886,306,1716) $DEVICE_ID=1003
MM6 36 2 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=336 $Y=1050  $PIN_XY=(366,1038,366,868),336,1050,(306,1038,306,868) $DEVICE_ID=1003
MM7 3 13 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=168 $Y=1704  $PIN_XY=(198,1886,198,1716),168,1704,(138,1886,138,1716) $DEVICE_ID=1003
MM8 4 2 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=168 $Y=1050  $PIN_XY=(198,1038,198,868),168,1050,(138,1038,138,868) $DEVICE_ID=1003
XX73A2B172333 13 3 34 35 38 41 inverter_column_decoder_write $T=-54 1394 0 0 $X=-54 $Y=1314
XX73A2B172334 2 4 34 36 38 42 inverter_column_decoder_write $T=-54 1360 1 0 $X=-54 $Y=660
XX73A2B172335_1 37 36 39 42 fill_sram_column_decoder_write $T=-30 70 0 0 $X=-54 $Y=6
XX73A2B172335_2 37 36 39 42 fill_sram_column_decoder_write $T=138 70 0 0 $X=114 $Y=6
XX73A2B172335_3 37 36 39 42 fill_sram_column_decoder_write $T=306 70 0 0 $X=282 $Y=6
XX73A2B172338 37 36 39 42 fill_sram_column_decoder_write $T=8202 70 0 0 $X=8178 $Y=6
XX73A2B172339_1 37 36 39 42 fill_sram_column_decoder_write $T=7194 70 0 0 $X=7170 $Y=6
XX73A2B172339_2 37 36 39 42 fill_sram_column_decoder_write $T=7362 70 0 0 $X=7338 $Y=6
XX73A2B172341_1 37 36 39 42 fill_sram_column_decoder_write $T=6186 70 0 0 $X=6162 $Y=6
XX73A2B172341_2 37 36 39 42 fill_sram_column_decoder_write $T=6354 70 0 0 $X=6330 $Y=6
XX73A2B172343_1 37 36 39 42 fill_sram_column_decoder_write $T=5178 70 0 0 $X=5154 $Y=6
XX73A2B172343_2 37 36 39 42 fill_sram_column_decoder_write $T=5346 70 0 0 $X=5322 $Y=6
XX73A2B172345_1 37 36 39 42 fill_sram_column_decoder_write $T=4170 70 0 0 $X=4146 $Y=6
XX73A2B172345_2 37 36 39 42 fill_sram_column_decoder_write $T=4338 70 0 0 $X=4314 $Y=6
XX73A2B172347_1 37 36 39 42 fill_sram_column_decoder_write $T=3162 70 0 0 $X=3138 $Y=6
XX73A2B172347_2 37 36 39 42 fill_sram_column_decoder_write $T=3330 70 0 0 $X=3306 $Y=6
XX73A2B172349_1 37 36 39 42 fill_sram_column_decoder_write $T=1146 70 0 0 $X=1122 $Y=6
XX73A2B172349_2 37 36 39 42 fill_sram_column_decoder_write $T=1314 70 0 0 $X=1290 $Y=6
XX73A2B172351_1 37 36 39 42 fill_sram_column_decoder_write $T=2154 70 0 0 $X=2130 $Y=6
XX73A2B172351_2 37 36 39 42 fill_sram_column_decoder_write $T=2322 70 0 0 $X=2298 $Y=6
XX73A2B172353 34 36 38 42 fill_sram_inverted $T=8202 1376 1 0 $X=8178 $Y=660
XX73A2B172354_1 34 36 38 42 fill_sram_inverted $T=6186 1376 1 0 $X=6162 $Y=660
XX73A2B172354_2 34 36 38 42 fill_sram_inverted $T=6354 1376 1 0 $X=6330 $Y=660
XX73A2B172356_1 34 36 38 42 fill_sram_inverted $T=4170 1376 1 0 $X=4146 $Y=660
XX73A2B172356_2 34 36 38 42 fill_sram_inverted $T=4338 1376 1 0 $X=4314 $Y=660
XX73A2B172358_1 34 36 38 42 fill_sram_inverted $T=2154 1376 1 0 $X=2130 $Y=660
XX73A2B172358_2 34 36 38 42 fill_sram_inverted $T=2322 1376 1 0 $X=2298 $Y=660
XX73A2B172360 2 6 4 14 15 37 36 39 42 column_decoder_write_cell $T=1458 0 0 0 $X=1458 $Y=6
XX73A2B172361 2 8 4 16 17 37 36 39 42 column_decoder_write_cell $T=3474 0 0 0 $X=3474 $Y=6
XX73A2B172362 2 5 4 18 19 37 36 39 42 column_decoder_write_cell $T=450 0 0 0 $X=450 $Y=6
XX73A2B172363 2 12 4 20 21 37 36 39 42 column_decoder_write_cell $T=7506 0 0 0 $X=7506 $Y=6
XX73A2B172364 2 11 4 22 23 37 36 39 42 column_decoder_write_cell $T=6498 0 0 0 $X=6498 $Y=6
XX73A2B172365 2 7 4 24 25 37 36 39 42 column_decoder_write_cell $T=2466 0 0 0 $X=2466 $Y=6
XX73A2B172366 2 10 4 26 27 37 36 39 42 column_decoder_write_cell $T=5490 0 0 0 $X=5490 $Y=6
XX73A2B172367 2 9 4 28 29 37 36 39 42 column_decoder_write_cell $T=4482 0 0 0 $X=4482 $Y=6
XX73A2B172368 34 35 38 41 fill_sram $T=8202 1378 0 0 $X=8178 $Y=1314
XX73A2B172369_1 34 35 38 41 fill_sram $T=4170 1378 0 0 $X=4146 $Y=1314
XX73A2B172369_2 34 35 38 41 fill_sram $T=4338 1378 0 0 $X=4314 $Y=1314
XX73A2B172371_1 34 35 38 41 fill_sram $T=2154 1378 0 0 $X=2130 $Y=1314
XX73A2B172371_2 34 35 38 41 fill_sram $T=2322 1378 0 0 $X=2298 $Y=1314
XX73A2B172373_1 34 35 38 41 fill_sram $T=6186 1378 0 0 $X=6162 $Y=1314
XX73A2B172373_2 34 35 38 41 fill_sram $T=6354 1378 0 0 $X=6330 $Y=1314
XX73A2B172375 30 3 11 12 34 35 36 38 40 41 42 write_buffer_cell $T=6216 2094 1 0 $X=6498 $Y=659
XX73A2B172376 31 3 9 10 34 35 36 38 40 41 42 write_buffer_cell $T=4200 2094 1 0 $X=4482 $Y=659
XX73A2B172377 32 3 7 8 34 35 36 38 40 41 42 write_buffer_cell $T=2184 2094 1 0 $X=2466 $Y=659
XX73A2B172378 33 3 5 6 34 35 36 38 40 41 42 write_buffer_cell $T=168 2094 1 0 $X=450 $Y=659
.ends column_decoder_write
.subckt VCELLR4 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 19 20 29 30 31
+	32 33 34 35 36 37 38 39 40 41 42
+	43 44 53 54 55 56 57 58 59 60 61
+	62 63 64 65 66 67 68 69 70 71 72
+	73 74 75 76 77 78 79
MM1 17 19 45 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3696 $Y=1454  $PIN_XY=3726,1452,3696,1454,3666,1452 $DEVICE_ID=1001
MM2 72 20 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3696 $Y=1160  $PIN_XY=3726,1162,3696,1160,3666,1162 $DEVICE_ID=1001
MM3 45 46 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3528 $Y=1634  $PIN_XY=3558,1452,3528,1634,3498,1452 $DEVICE_ID=1001
MM4 21 22 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3528 $Y=980  $PIN_XY=3558,1162,3528,980,3498,1162 $DEVICE_ID=1001
MM5 55 45 46 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3360 $Y=1634  $PIN_XY=3390,1452,3360,1634,3330,1452 $DEVICE_ID=1001
MM6 55 21 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3360 $Y=980  $PIN_XY=3390,1162,3360,980,3330,1162 $DEVICE_ID=1001
MM7 46 19 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=1454  $PIN_XY=3222,1452,3192,1454,3162,1452 $DEVICE_ID=1001
MM8 22 20 71 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=1160  $PIN_XY=3222,1162,3192,1160,3162,1162 $DEVICE_ID=1001
MM9 13 19 47 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2688 $Y=1454  $PIN_XY=2718,1452,2688,1454,2658,1452 $DEVICE_ID=1001
MM10 69 20 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2688 $Y=1160  $PIN_XY=2718,1162,2688,1160,2658,1162 $DEVICE_ID=1001
MM11 47 48 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2520 $Y=1634  $PIN_XY=2550,1452,2520,1634,2490,1452 $DEVICE_ID=1001
MM12 23 24 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2520 $Y=980  $PIN_XY=2550,1162,2520,980,2490,1162 $DEVICE_ID=1001
MM13 55 47 48 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2352 $Y=1634  $PIN_XY=2382,1452,2352,1634,2322,1452 $DEVICE_ID=1001
MM14 55 23 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2352 $Y=980  $PIN_XY=2382,1162,2352,980,2322,1162 $DEVICE_ID=1001
MM15 48 19 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2184 $Y=1454  $PIN_XY=2214,1452,2184,1454,2154,1452 $DEVICE_ID=1001
MM16 24 20 68 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2184 $Y=1160  $PIN_XY=2214,1162,2184,1160,2154,1162 $DEVICE_ID=1001
MM17 9 19 49 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1680 $Y=1454  $PIN_XY=1710,1452,1680,1454,1650,1452 $DEVICE_ID=1001
MM18 67 20 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1680 $Y=1160  $PIN_XY=1710,1162,1680,1160,1650,1162 $DEVICE_ID=1001
MM19 49 50 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1512 $Y=1634  $PIN_XY=1542,1452,1512,1634,1482,1452 $DEVICE_ID=1001
MM20 25 26 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1512 $Y=980  $PIN_XY=1542,1162,1512,980,1482,1162 $DEVICE_ID=1001
MM21 55 49 50 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1344 $Y=1634  $PIN_XY=1374,1452,1344,1634,1314,1452 $DEVICE_ID=1001
MM22 55 25 26 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1344 $Y=980  $PIN_XY=1374,1162,1344,980,1314,1162 $DEVICE_ID=1001
MM23 50 19 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1176 $Y=1454  $PIN_XY=1206,1452,1176,1454,1146,1452 $DEVICE_ID=1001
MM24 26 20 70 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1176 $Y=1160  $PIN_XY=1206,1162,1176,1160,1146,1162 $DEVICE_ID=1001
MM25 5 19 51 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=672 $Y=1454  $PIN_XY=702,1452,672,1454,642,1452 $DEVICE_ID=1001
MM26 66 20 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=672 $Y=1160  $PIN_XY=702,1162,672,1160,642,1162 $DEVICE_ID=1001
MM27 51 52 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=504 $Y=1634  $PIN_XY=534,1452,504,1634,474,1452 $DEVICE_ID=1001
MM28 27 28 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=504 $Y=980  $PIN_XY=534,1162,504,980,474,1162 $DEVICE_ID=1001
MM29 55 51 52 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=1634  $PIN_XY=366,1452,336,1634,306,1452 $DEVICE_ID=1001
MM30 55 27 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=980  $PIN_XY=366,1162,336,980,306,1162 $DEVICE_ID=1001
MM31 52 19 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=1454  $PIN_XY=198,1452,168,1454,138,1452 $DEVICE_ID=1001
MM32 28 20 65 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=1160  $PIN_XY=198,1162,168,1160,138,1162 $DEVICE_ID=1001
MM33 29 30 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3528 $Y=2288  $PIN_XY=(3558,2276,3558,2106),3528,2288,(3498,2276,3498,2106) $DEVICE_ID=1003
MM34 45 46 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3528 $Y=1634  $PIN_XY=(3558,1816,3558,1646),3528,1634,(3498,1816,3498,1646) $DEVICE_ID=1003
MM35 21 22 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3528 $Y=980  $PIN_XY=(3558,968,3558,798),3528,980,(3498,968,3498,798) $DEVICE_ID=1003
MM36 37 38 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3528 $Y=326  $PIN_XY=(3558,508,3558,338),3528,326,(3498,508,3498,338) $DEVICE_ID=1003
MM37 54 29 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3360 $Y=2288  $PIN_XY=(3390,2276,3390,2106),3360,2288,(3330,2276,3330,2106) $DEVICE_ID=1003
MM38 54 45 46 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3360 $Y=1634  $PIN_XY=(3390,1816,3390,1646),3360,1634,(3330,1816,3330,1646) $DEVICE_ID=1003
MM39 53 21 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3360 $Y=980  $PIN_XY=(3390,968,3390,798),3360,980,(3330,968,3330,798) $DEVICE_ID=1003
MM40 53 37 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3360 $Y=326  $PIN_XY=(3390,508,3390,338),3360,326,(3330,508,3330,338) $DEVICE_ID=1003
MM41 31 32 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=2520 $Y=2288  $PIN_XY=(2550,2276,2550,2106),2520,2288,(2490,2276,2490,2106) $DEVICE_ID=1003
MM42 47 48 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=2520 $Y=1634  $PIN_XY=(2550,1816,2550,1646),2520,1634,(2490,1816,2490,1646) $DEVICE_ID=1003
MM43 23 24 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=2520 $Y=980  $PIN_XY=(2550,968,2550,798),2520,980,(2490,968,2490,798) $DEVICE_ID=1003
MM44 39 40 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=2520 $Y=326  $PIN_XY=(2550,508,2550,338),2520,326,(2490,508,2490,338) $DEVICE_ID=1003
MM45 54 31 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=2352 $Y=2288  $PIN_XY=(2382,2276,2382,2106),2352,2288,(2322,2276,2322,2106) $DEVICE_ID=1003
MM46 54 47 48 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=2352 $Y=1634  $PIN_XY=(2382,1816,2382,1646),2352,1634,(2322,1816,2322,1646) $DEVICE_ID=1003
MM47 53 23 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=2352 $Y=980  $PIN_XY=(2382,968,2382,798),2352,980,(2322,968,2322,798) $DEVICE_ID=1003
MM48 53 39 40 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=2352 $Y=326  $PIN_XY=(2382,508,2382,338),2352,326,(2322,508,2322,338) $DEVICE_ID=1003
MM49 33 34 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=1512 $Y=2288  $PIN_XY=(1542,2276,1542,2106),1512,2288,(1482,2276,1482,2106) $DEVICE_ID=1003
MM50 49 50 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=1512 $Y=1634  $PIN_XY=(1542,1816,1542,1646),1512,1634,(1482,1816,1482,1646) $DEVICE_ID=1003
MM51 25 26 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=1512 $Y=980  $PIN_XY=(1542,968,1542,798),1512,980,(1482,968,1482,798) $DEVICE_ID=1003
MM52 41 42 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=1512 $Y=326  $PIN_XY=(1542,508,1542,338),1512,326,(1482,508,1482,338) $DEVICE_ID=1003
MM53 54 33 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=1344 $Y=2288  $PIN_XY=(1374,2276,1374,2106),1344,2288,(1314,2276,1314,2106) $DEVICE_ID=1003
MM54 54 49 50 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=1344 $Y=1634  $PIN_XY=(1374,1816,1374,1646),1344,1634,(1314,1816,1314,1646) $DEVICE_ID=1003
MM55 53 25 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=1344 $Y=980  $PIN_XY=(1374,968,1374,798),1344,980,(1314,968,1314,798) $DEVICE_ID=1003
MM56 53 41 42 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=1344 $Y=326  $PIN_XY=(1374,508,1374,338),1344,326,(1314,508,1314,338) $DEVICE_ID=1003
MM57 35 36 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=504 $Y=2288  $PIN_XY=(534,2276,534,2106),504,2288,(474,2276,474,2106) $DEVICE_ID=1003
MM58 51 52 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=504 $Y=1634  $PIN_XY=(534,1816,534,1646),504,1634,(474,1816,474,1646) $DEVICE_ID=1003
MM59 27 28 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=504 $Y=980  $PIN_XY=(534,968,534,798),504,980,(474,968,474,798) $DEVICE_ID=1003
MM60 43 44 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=504 $Y=326  $PIN_XY=(534,508,534,338),504,326,(474,508,474,338) $DEVICE_ID=1003
MM61 54 35 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=336 $Y=2288  $PIN_XY=(366,2276,366,2106),336,2288,(306,2276,306,2106) $DEVICE_ID=1003
MM62 54 51 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=336 $Y=1634  $PIN_XY=(366,1816,366,1646),336,1634,(306,1816,306,1646) $DEVICE_ID=1003
MM63 53 27 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=336 $Y=980  $PIN_XY=(366,968,366,798),336,980,(306,968,306,798) $DEVICE_ID=1003
MM64 53 43 44 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=336 $Y=326  $PIN_XY=(366,508,366,338),336,326,(306,508,306,338) $DEVICE_ID=1003
XX73A2B172452 65 66 70 67 68 69 71 72 20 55 53 
+	21 22 23 24 25 26 27 28 75 77 sram_array_1r_4c $T=0 1306 1 0 $X=-54 $Y=590
XX73A2B172453 57 58 62 59 60 61 63 64 73 74 54 
+	29 30 31 32 33 34 35 36 79 78 sram_array_1r_4c $T=0 2614 1 0 $X=-54 $Y=1898
XX73A2B172454 14 18 16 38 37 53 56 76 77 sram_6T_1finger_inverted $T=3024 16 0 0 $X=2970 $Y=-64
XX73A2B172455 10 18 12 40 39 53 56 76 77 sram_6T_1finger_inverted $T=2016 16 0 0 $X=1962 $Y=-64
XX73A2B172456 6 18 8 42 41 53 56 76 77 sram_6T_1finger_inverted $T=1008 16 0 0 $X=954 $Y=-64
XX73A2B172457 2 18 4 44 43 53 56 76 77 sram_6T_1finger_inverted $T=0 16 0 0 $X=-54 $Y=-64
XX73A2B172458 15 19 17 46 45 54 55 75 78 sram_6T_1finger_inverted $T=3024 1324 0 0 $X=2970 $Y=1244
XX73A2B172459 11 19 13 48 47 54 55 75 78 sram_6T_1finger_inverted $T=2016 1324 0 0 $X=1962 $Y=1244
XX73A2B172460 7 19 9 50 49 54 55 75 78 sram_6T_1finger_inverted $T=1008 1324 0 0 $X=954 $Y=1244
XX73A2B172461 3 19 5 52 51 54 55 75 78 sram_6T_1finger_inverted $T=0 1324 0 0 $X=-54 $Y=1244
XX73A2B172462 56 53 76 77 fill_sram_inverted $T=2826 0 0 0 $X=2802 $Y=-64
XX73A2B172463 56 53 76 77 fill_sram_inverted $T=1818 0 0 0 $X=1794 $Y=-64
XX73A2B172464 56 53 76 77 fill_sram_inverted $T=810 0 0 0 $X=786 $Y=-64
XX73A2B172465 55 54 75 78 fill_sram_inverted $T=2826 1308 0 0 $X=2802 $Y=1244
XX73A2B172466 55 54 75 78 fill_sram_inverted $T=1818 1308 0 0 $X=1794 $Y=1244
XX73A2B172467 55 54 75 78 fill_sram_inverted $T=810 1308 0 0 $X=786 $Y=1244
.ends VCELLR4

* Hierarchy Level 1
.subckt sram_array_16r_8c 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 23
+	24 25 26 27 28 29 30 31 32 33 130
+	131 132 133 134 135 136 137 138 139 140 141
+	142 143 144 145 146 147 148 149 150 151 152
+	153 154 155 156 157 158 159 160 161 162 163
+	164 165 166 167 168 169 170 171 172 173 174
+	175 176 177 178 179 180 181 182 183 184 185
+	186 187 188 189 190 191 192 193 194 195
MM1 17 33 122 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=7994  $PIN_XY=7758,7992,7728,7994,7698,7992 $DEVICE_ID=1001
MM2 17 26 114 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=7700  $PIN_XY=7758,7702,7728,7700,7698,7702 $DEVICE_ID=1001
MM3 17 29 106 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=5378  $PIN_XY=7758,5376,7728,5378,7698,5376 $DEVICE_ID=1001
MM4 17 22 98 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=5084  $PIN_XY=7758,5086,7728,5084,7698,5086 $DEVICE_ID=1001
MM5 122 123 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7560 $Y=8174  $PIN_XY=7590,7992,7560,8174,7530,7992 $DEVICE_ID=1001
MM6 114 115 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7560 $Y=7520  $PIN_XY=7590,7702,7560,7520,7530,7702 $DEVICE_ID=1001
MM7 106 107 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7560 $Y=5558  $PIN_XY=7590,5376,7560,5558,7530,5376 $DEVICE_ID=1001
MM8 98 99 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7560 $Y=4904  $PIN_XY=7590,5086,7560,4904,7530,5086 $DEVICE_ID=1001
MM9 133 122 123 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7392 $Y=8174  $PIN_XY=7422,7992,7392,8174,7362,7992 $DEVICE_ID=1001
MM10 133 114 115 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7392 $Y=7520  $PIN_XY=7422,7702,7392,7520,7362,7702 $DEVICE_ID=1001
MM11 140 106 107 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7392 $Y=5558  $PIN_XY=7422,5376,7392,5558,7362,5376 $DEVICE_ID=1001
MM12 140 98 99 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7392 $Y=4904  $PIN_XY=7422,5086,7392,4904,7362,5086 $DEVICE_ID=1001
MM13 123 33 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7224 $Y=7994  $PIN_XY=7254,7992,7224,7994,7194,7992 $DEVICE_ID=1001
MM14 115 26 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7224 $Y=7700  $PIN_XY=7254,7702,7224,7700,7194,7702 $DEVICE_ID=1001
MM15 107 29 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7224 $Y=5378  $PIN_XY=7254,5376,7224,5378,7194,5376 $DEVICE_ID=1001
MM16 99 22 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7224 $Y=5084  $PIN_XY=7254,5086,7224,5084,7194,5086 $DEVICE_ID=1001
MM17 15 33 124 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6720 $Y=7994  $PIN_XY=6750,7992,6720,7994,6690,7992 $DEVICE_ID=1001
MM18 15 26 116 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6720 $Y=7700  $PIN_XY=6750,7702,6720,7700,6690,7702 $DEVICE_ID=1001
MM19 15 29 108 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6720 $Y=5378  $PIN_XY=6750,5376,6720,5378,6690,5376 $DEVICE_ID=1001
MM20 15 22 100 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6720 $Y=5084  $PIN_XY=6750,5086,6720,5084,6690,5086 $DEVICE_ID=1001
MM21 124 125 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6552 $Y=8174  $PIN_XY=6582,7992,6552,8174,6522,7992 $DEVICE_ID=1001
MM22 116 117 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6552 $Y=7520  $PIN_XY=6582,7702,6552,7520,6522,7702 $DEVICE_ID=1001
MM23 108 109 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6552 $Y=5558  $PIN_XY=6582,5376,6552,5558,6522,5376 $DEVICE_ID=1001
MM24 100 101 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6552 $Y=4904  $PIN_XY=6582,5086,6552,4904,6522,5086 $DEVICE_ID=1001
MM25 133 124 125 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6384 $Y=8174  $PIN_XY=6414,7992,6384,8174,6354,7992 $DEVICE_ID=1001
MM26 133 116 117 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6384 $Y=7520  $PIN_XY=6414,7702,6384,7520,6354,7702 $DEVICE_ID=1001
MM27 140 108 109 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6384 $Y=5558  $PIN_XY=6414,5376,6384,5558,6354,5376 $DEVICE_ID=1001
MM28 140 100 101 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6384 $Y=4904  $PIN_XY=6414,5086,6384,4904,6354,5086 $DEVICE_ID=1001
MM29 125 33 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6216 $Y=7994  $PIN_XY=6246,7992,6216,7994,6186,7992 $DEVICE_ID=1001
MM30 117 26 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6216 $Y=7700  $PIN_XY=6246,7702,6216,7700,6186,7702 $DEVICE_ID=1001
MM31 109 29 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6216 $Y=5378  $PIN_XY=6246,5376,6216,5378,6186,5376 $DEVICE_ID=1001
MM32 101 22 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6216 $Y=5084  $PIN_XY=6246,5086,6216,5084,6186,5086 $DEVICE_ID=1001
MM33 13 33 126 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5712 $Y=7994  $PIN_XY=5742,7992,5712,7994,5682,7992 $DEVICE_ID=1001
MM34 13 26 118 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5712 $Y=7700  $PIN_XY=5742,7702,5712,7700,5682,7702 $DEVICE_ID=1001
MM35 13 29 110 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5712 $Y=5378  $PIN_XY=5742,5376,5712,5378,5682,5376 $DEVICE_ID=1001
MM36 13 22 102 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5712 $Y=5084  $PIN_XY=5742,5086,5712,5084,5682,5086 $DEVICE_ID=1001
MM37 126 127 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5544 $Y=8174  $PIN_XY=5574,7992,5544,8174,5514,7992 $DEVICE_ID=1001
MM38 118 119 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5544 $Y=7520  $PIN_XY=5574,7702,5544,7520,5514,7702 $DEVICE_ID=1001
MM39 110 111 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5544 $Y=5558  $PIN_XY=5574,5376,5544,5558,5514,5376 $DEVICE_ID=1001
MM40 102 103 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5544 $Y=4904  $PIN_XY=5574,5086,5544,4904,5514,5086 $DEVICE_ID=1001
MM41 133 126 127 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5376 $Y=8174  $PIN_XY=5406,7992,5376,8174,5346,7992 $DEVICE_ID=1001
MM42 133 118 119 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5376 $Y=7520  $PIN_XY=5406,7702,5376,7520,5346,7702 $DEVICE_ID=1001
MM43 140 110 111 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5376 $Y=5558  $PIN_XY=5406,5376,5376,5558,5346,5376 $DEVICE_ID=1001
MM44 140 102 103 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5376 $Y=4904  $PIN_XY=5406,5086,5376,4904,5346,5086 $DEVICE_ID=1001
MM45 127 33 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5208 $Y=7994  $PIN_XY=5238,7992,5208,7994,5178,7992 $DEVICE_ID=1001
MM46 119 26 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5208 $Y=7700  $PIN_XY=5238,7702,5208,7700,5178,7702 $DEVICE_ID=1001
MM47 111 29 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5208 $Y=5378  $PIN_XY=5238,5376,5208,5378,5178,5376 $DEVICE_ID=1001
MM48 103 22 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5208 $Y=5084  $PIN_XY=5238,5086,5208,5084,5178,5086 $DEVICE_ID=1001
MM49 11 33 128 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4704 $Y=7994  $PIN_XY=4734,7992,4704,7994,4674,7992 $DEVICE_ID=1001
MM50 11 26 120 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4704 $Y=7700  $PIN_XY=4734,7702,4704,7700,4674,7702 $DEVICE_ID=1001
MM51 11 29 112 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4704 $Y=5378  $PIN_XY=4734,5376,4704,5378,4674,5376 $DEVICE_ID=1001
MM52 11 22 104 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4704 $Y=5084  $PIN_XY=4734,5086,4704,5084,4674,5086 $DEVICE_ID=1001
MM53 128 129 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4536 $Y=8174  $PIN_XY=4566,7992,4536,8174,4506,7992 $DEVICE_ID=1001
MM54 120 121 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4536 $Y=7520  $PIN_XY=4566,7702,4536,7520,4506,7702 $DEVICE_ID=1001
MM55 112 113 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4536 $Y=5558  $PIN_XY=4566,5376,4536,5558,4506,5376 $DEVICE_ID=1001
MM56 104 105 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4536 $Y=4904  $PIN_XY=4566,5086,4536,4904,4506,5086 $DEVICE_ID=1001
MM57 133 128 129 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4368 $Y=8174  $PIN_XY=4398,7992,4368,8174,4338,7992 $DEVICE_ID=1001
MM58 133 120 121 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4368 $Y=7520  $PIN_XY=4398,7702,4368,7520,4338,7702 $DEVICE_ID=1001
MM59 140 112 113 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4368 $Y=5558  $PIN_XY=4398,5376,4368,5558,4338,5376 $DEVICE_ID=1001
MM60 140 104 105 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4368 $Y=4904  $PIN_XY=4398,5086,4368,4904,4338,5086 $DEVICE_ID=1001
MM61 129 33 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=7994  $PIN_XY=4230,7992,4200,7994,4170,7992 $DEVICE_ID=1001
MM62 121 26 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=7700  $PIN_XY=4230,7702,4200,7700,4170,7702 $DEVICE_ID=1001
MM63 113 29 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=5378  $PIN_XY=4230,5376,4200,5378,4170,5376 $DEVICE_ID=1001
MM64 105 22 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=5084  $PIN_XY=4230,5086,4200,5084,4170,5086 $DEVICE_ID=1001
MM65 9 33 74 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3696 $Y=7994  $PIN_XY=3726,7992,3696,7994,3666,7992 $DEVICE_ID=1001
MM66 9 26 66 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3696 $Y=7700  $PIN_XY=3726,7702,3696,7700,3666,7702 $DEVICE_ID=1001
MM67 9 29 58 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3696 $Y=5378  $PIN_XY=3726,5376,3696,5378,3666,5376 $DEVICE_ID=1001
MM68 9 22 50 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3696 $Y=5084  $PIN_XY=3726,5086,3696,5084,3666,5086 $DEVICE_ID=1001
MM69 74 75 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3528 $Y=8174  $PIN_XY=3558,7992,3528,8174,3498,7992 $DEVICE_ID=1001
MM70 66 67 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3528 $Y=7520  $PIN_XY=3558,7702,3528,7520,3498,7702 $DEVICE_ID=1001
MM71 58 59 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3528 $Y=5558  $PIN_XY=3558,5376,3528,5558,3498,5376 $DEVICE_ID=1001
MM72 50 51 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3528 $Y=4904  $PIN_XY=3558,5086,3528,4904,3498,5086 $DEVICE_ID=1001
MM73 133 74 75 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3360 $Y=8174  $PIN_XY=3390,7992,3360,8174,3330,7992 $DEVICE_ID=1001
MM74 133 66 67 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3360 $Y=7520  $PIN_XY=3390,7702,3360,7520,3330,7702 $DEVICE_ID=1001
MM75 140 58 59 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3360 $Y=5558  $PIN_XY=3390,5376,3360,5558,3330,5376 $DEVICE_ID=1001
MM76 140 50 51 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3360 $Y=4904  $PIN_XY=3390,5086,3360,4904,3330,5086 $DEVICE_ID=1001
MM77 75 33 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=7994  $PIN_XY=3222,7992,3192,7994,3162,7992 $DEVICE_ID=1001
MM78 67 26 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=7700  $PIN_XY=3222,7702,3192,7700,3162,7702 $DEVICE_ID=1001
MM79 59 29 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=5378  $PIN_XY=3222,5376,3192,5378,3162,5376 $DEVICE_ID=1001
MM80 51 22 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=5084  $PIN_XY=3222,5086,3192,5084,3162,5086 $DEVICE_ID=1001
MM81 7 33 76 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2688 $Y=7994  $PIN_XY=2718,7992,2688,7994,2658,7992 $DEVICE_ID=1001
MM82 7 26 68 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2688 $Y=7700  $PIN_XY=2718,7702,2688,7700,2658,7702 $DEVICE_ID=1001
MM83 7 29 60 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2688 $Y=5378  $PIN_XY=2718,5376,2688,5378,2658,5376 $DEVICE_ID=1001
MM84 7 22 52 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2688 $Y=5084  $PIN_XY=2718,5086,2688,5084,2658,5086 $DEVICE_ID=1001
MM85 76 77 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2520 $Y=8174  $PIN_XY=2550,7992,2520,8174,2490,7992 $DEVICE_ID=1001
MM86 68 69 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2520 $Y=7520  $PIN_XY=2550,7702,2520,7520,2490,7702 $DEVICE_ID=1001
MM87 60 61 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2520 $Y=5558  $PIN_XY=2550,5376,2520,5558,2490,5376 $DEVICE_ID=1001
MM88 52 53 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2520 $Y=4904  $PIN_XY=2550,5086,2520,4904,2490,5086 $DEVICE_ID=1001
MM89 133 76 77 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2352 $Y=8174  $PIN_XY=2382,7992,2352,8174,2322,7992 $DEVICE_ID=1001
MM90 133 68 69 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2352 $Y=7520  $PIN_XY=2382,7702,2352,7520,2322,7702 $DEVICE_ID=1001
MM91 140 60 61 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2352 $Y=5558  $PIN_XY=2382,5376,2352,5558,2322,5376 $DEVICE_ID=1001
MM92 140 52 53 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2352 $Y=4904  $PIN_XY=2382,5086,2352,4904,2322,5086 $DEVICE_ID=1001
MM93 77 33 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2184 $Y=7994  $PIN_XY=2214,7992,2184,7994,2154,7992 $DEVICE_ID=1001
MM94 69 26 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2184 $Y=7700  $PIN_XY=2214,7702,2184,7700,2154,7702 $DEVICE_ID=1001
MM95 61 29 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2184 $Y=5378  $PIN_XY=2214,5376,2184,5378,2154,5376 $DEVICE_ID=1001
MM96 53 22 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2184 $Y=5084  $PIN_XY=2214,5086,2184,5084,2154,5086 $DEVICE_ID=1001
MM97 5 33 78 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1680 $Y=7994  $PIN_XY=1710,7992,1680,7994,1650,7992 $DEVICE_ID=1001
MM98 5 26 70 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1680 $Y=7700  $PIN_XY=1710,7702,1680,7700,1650,7702 $DEVICE_ID=1001
MM99 5 29 62 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1680 $Y=5378  $PIN_XY=1710,5376,1680,5378,1650,5376 $DEVICE_ID=1001
MM100 5 22 54 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1680 $Y=5084  $PIN_XY=1710,5086,1680,5084,1650,5086 $DEVICE_ID=1001
MM101 78 79 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1512 $Y=8174  $PIN_XY=1542,7992,1512,8174,1482,7992 $DEVICE_ID=1001
MM102 70 71 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1512 $Y=7520  $PIN_XY=1542,7702,1512,7520,1482,7702 $DEVICE_ID=1001
MM103 62 63 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1512 $Y=5558  $PIN_XY=1542,5376,1512,5558,1482,5376 $DEVICE_ID=1001
MM104 54 55 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1512 $Y=4904  $PIN_XY=1542,5086,1512,4904,1482,5086 $DEVICE_ID=1001
MM105 133 78 79 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1344 $Y=8174  $PIN_XY=1374,7992,1344,8174,1314,7992 $DEVICE_ID=1001
MM106 133 70 71 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1344 $Y=7520  $PIN_XY=1374,7702,1344,7520,1314,7702 $DEVICE_ID=1001
MM107 140 62 63 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1344 $Y=5558  $PIN_XY=1374,5376,1344,5558,1314,5376 $DEVICE_ID=1001
MM108 140 54 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1344 $Y=4904  $PIN_XY=1374,5086,1344,4904,1314,5086 $DEVICE_ID=1001
MM109 79 33 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1176 $Y=7994  $PIN_XY=1206,7992,1176,7994,1146,7992 $DEVICE_ID=1001
MM110 71 26 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1176 $Y=7700  $PIN_XY=1206,7702,1176,7700,1146,7702 $DEVICE_ID=1001
MM111 63 29 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1176 $Y=5378  $PIN_XY=1206,5376,1176,5378,1146,5376 $DEVICE_ID=1001
MM112 55 22 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1176 $Y=5084  $PIN_XY=1206,5086,1176,5084,1146,5086 $DEVICE_ID=1001
MM113 3 33 80 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=672 $Y=7994  $PIN_XY=702,7992,672,7994,642,7992 $DEVICE_ID=1001
MM114 3 26 72 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=672 $Y=7700  $PIN_XY=702,7702,672,7700,642,7702 $DEVICE_ID=1001
MM115 3 29 64 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=672 $Y=5378  $PIN_XY=702,5376,672,5378,642,5376 $DEVICE_ID=1001
MM116 3 22 56 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=672 $Y=5084  $PIN_XY=702,5086,672,5084,642,5086 $DEVICE_ID=1001
MM117 80 81 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=504 $Y=8174  $PIN_XY=534,7992,504,8174,474,7992 $DEVICE_ID=1001
MM118 72 73 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=504 $Y=7520  $PIN_XY=534,7702,504,7520,474,7702 $DEVICE_ID=1001
MM119 64 65 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=504 $Y=5558  $PIN_XY=534,5376,504,5558,474,5376 $DEVICE_ID=1001
MM120 56 57 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=504 $Y=4904  $PIN_XY=534,5086,504,4904,474,5086 $DEVICE_ID=1001
MM121 133 80 81 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=8174  $PIN_XY=366,7992,336,8174,306,7992 $DEVICE_ID=1001
MM122 133 72 73 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=7520  $PIN_XY=366,7702,336,7520,306,7702 $DEVICE_ID=1001
MM123 140 64 65 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=5558  $PIN_XY=366,5376,336,5558,306,5376 $DEVICE_ID=1001
MM124 140 56 57 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=4904  $PIN_XY=366,5086,336,4904,306,5086 $DEVICE_ID=1001
MM125 81 33 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=7994  $PIN_XY=198,7992,168,7994,138,7992 $DEVICE_ID=1001
MM126 73 26 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=7700  $PIN_XY=198,7702,168,7700,138,7702 $DEVICE_ID=1001
MM127 65 29 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=5378  $PIN_XY=198,5376,168,5378,138,5376 $DEVICE_ID=1001
MM128 57 22 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=5084  $PIN_XY=198,5086,168,5084,138,5086 $DEVICE_ID=1001
MM129 17 25 90 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=2762  $PIN_XY=7758,2760,7728,2762,7698,2760 $DEVICE_ID=1001
MM130 17 18 82 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=2468  $PIN_XY=7758,2470,7728,2468,7698,2470 $DEVICE_ID=1001
MM131 90 91 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7560 $Y=2942  $PIN_XY=7590,2760,7560,2942,7530,2760 $DEVICE_ID=1001
MM132 82 83 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7560 $Y=2288  $PIN_XY=7590,2470,7560,2288,7530,2470 $DEVICE_ID=1001
MM133 142 90 91 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7392 $Y=2942  $PIN_XY=7422,2760,7392,2942,7362,2760 $DEVICE_ID=1001
MM134 142 82 83 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7392 $Y=2288  $PIN_XY=7422,2470,7392,2288,7362,2470 $DEVICE_ID=1001
MM135 91 25 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7224 $Y=2762  $PIN_XY=7254,2760,7224,2762,7194,2760 $DEVICE_ID=1001
MM136 83 18 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7224 $Y=2468  $PIN_XY=7254,2470,7224,2468,7194,2470 $DEVICE_ID=1001
MM137 15 25 92 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6720 $Y=2762  $PIN_XY=6750,2760,6720,2762,6690,2760 $DEVICE_ID=1001
MM138 15 18 84 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6720 $Y=2468  $PIN_XY=6750,2470,6720,2468,6690,2470 $DEVICE_ID=1001
MM139 92 93 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6552 $Y=2942  $PIN_XY=6582,2760,6552,2942,6522,2760 $DEVICE_ID=1001
MM140 84 85 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6552 $Y=2288  $PIN_XY=6582,2470,6552,2288,6522,2470 $DEVICE_ID=1001
MM141 142 92 93 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6384 $Y=2942  $PIN_XY=6414,2760,6384,2942,6354,2760 $DEVICE_ID=1001
MM142 142 84 85 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6384 $Y=2288  $PIN_XY=6414,2470,6384,2288,6354,2470 $DEVICE_ID=1001
MM143 93 25 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6216 $Y=2762  $PIN_XY=6246,2760,6216,2762,6186,2760 $DEVICE_ID=1001
MM144 85 18 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6216 $Y=2468  $PIN_XY=6246,2470,6216,2468,6186,2470 $DEVICE_ID=1001
MM145 13 25 94 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5712 $Y=2762  $PIN_XY=5742,2760,5712,2762,5682,2760 $DEVICE_ID=1001
MM146 13 18 86 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5712 $Y=2468  $PIN_XY=5742,2470,5712,2468,5682,2470 $DEVICE_ID=1001
MM147 94 95 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5544 $Y=2942  $PIN_XY=5574,2760,5544,2942,5514,2760 $DEVICE_ID=1001
MM148 86 87 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5544 $Y=2288  $PIN_XY=5574,2470,5544,2288,5514,2470 $DEVICE_ID=1001
MM149 142 94 95 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5376 $Y=2942  $PIN_XY=5406,2760,5376,2942,5346,2760 $DEVICE_ID=1001
MM150 142 86 87 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5376 $Y=2288  $PIN_XY=5406,2470,5376,2288,5346,2470 $DEVICE_ID=1001
MM151 95 25 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5208 $Y=2762  $PIN_XY=5238,2760,5208,2762,5178,2760 $DEVICE_ID=1001
MM152 87 18 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5208 $Y=2468  $PIN_XY=5238,2470,5208,2468,5178,2470 $DEVICE_ID=1001
MM153 11 25 96 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4704 $Y=2762  $PIN_XY=4734,2760,4704,2762,4674,2760 $DEVICE_ID=1001
MM154 11 18 88 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4704 $Y=2468  $PIN_XY=4734,2470,4704,2468,4674,2470 $DEVICE_ID=1001
MM155 96 97 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4536 $Y=2942  $PIN_XY=4566,2760,4536,2942,4506,2760 $DEVICE_ID=1001
MM156 88 89 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4536 $Y=2288  $PIN_XY=4566,2470,4536,2288,4506,2470 $DEVICE_ID=1001
MM157 142 96 97 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4368 $Y=2942  $PIN_XY=4398,2760,4368,2942,4338,2760 $DEVICE_ID=1001
MM158 142 88 89 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4368 $Y=2288  $PIN_XY=4398,2470,4368,2288,4338,2470 $DEVICE_ID=1001
MM159 97 25 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=2762  $PIN_XY=4230,2760,4200,2762,4170,2760 $DEVICE_ID=1001
MM160 89 18 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=2468  $PIN_XY=4230,2470,4200,2468,4170,2470 $DEVICE_ID=1001
MM161 9 25 42 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3696 $Y=2762  $PIN_XY=3726,2760,3696,2762,3666,2760 $DEVICE_ID=1001
MM162 9 18 34 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3696 $Y=2468  $PIN_XY=3726,2470,3696,2468,3666,2470 $DEVICE_ID=1001
MM163 42 43 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3528 $Y=2942  $PIN_XY=3558,2760,3528,2942,3498,2760 $DEVICE_ID=1001
MM164 34 35 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3528 $Y=2288  $PIN_XY=3558,2470,3528,2288,3498,2470 $DEVICE_ID=1001
MM165 142 42 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3360 $Y=2942  $PIN_XY=3390,2760,3360,2942,3330,2760 $DEVICE_ID=1001
MM166 142 34 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3360 $Y=2288  $PIN_XY=3390,2470,3360,2288,3330,2470 $DEVICE_ID=1001
MM167 43 25 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=2762  $PIN_XY=3222,2760,3192,2762,3162,2760 $DEVICE_ID=1001
MM168 35 18 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=2468  $PIN_XY=3222,2470,3192,2468,3162,2470 $DEVICE_ID=1001
MM169 7 25 44 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2688 $Y=2762  $PIN_XY=2718,2760,2688,2762,2658,2760 $DEVICE_ID=1001
MM170 7 18 36 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2688 $Y=2468  $PIN_XY=2718,2470,2688,2468,2658,2470 $DEVICE_ID=1001
MM171 44 45 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2520 $Y=2942  $PIN_XY=2550,2760,2520,2942,2490,2760 $DEVICE_ID=1001
MM172 36 37 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2520 $Y=2288  $PIN_XY=2550,2470,2520,2288,2490,2470 $DEVICE_ID=1001
MM173 142 44 45 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2352 $Y=2942  $PIN_XY=2382,2760,2352,2942,2322,2760 $DEVICE_ID=1001
MM174 142 36 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2352 $Y=2288  $PIN_XY=2382,2470,2352,2288,2322,2470 $DEVICE_ID=1001
MM175 45 25 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2184 $Y=2762  $PIN_XY=2214,2760,2184,2762,2154,2760 $DEVICE_ID=1001
MM176 37 18 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2184 $Y=2468  $PIN_XY=2214,2470,2184,2468,2154,2470 $DEVICE_ID=1001
MM177 5 25 46 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1680 $Y=2762  $PIN_XY=1710,2760,1680,2762,1650,2760 $DEVICE_ID=1001
MM178 5 18 38 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1680 $Y=2468  $PIN_XY=1710,2470,1680,2468,1650,2470 $DEVICE_ID=1001
MM179 46 47 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1512 $Y=2942  $PIN_XY=1542,2760,1512,2942,1482,2760 $DEVICE_ID=1001
MM180 38 39 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1512 $Y=2288  $PIN_XY=1542,2470,1512,2288,1482,2470 $DEVICE_ID=1001
MM181 142 46 47 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1344 $Y=2942  $PIN_XY=1374,2760,1344,2942,1314,2760 $DEVICE_ID=1001
MM182 142 38 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1344 $Y=2288  $PIN_XY=1374,2470,1344,2288,1314,2470 $DEVICE_ID=1001
MM183 47 25 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1176 $Y=2762  $PIN_XY=1206,2760,1176,2762,1146,2760 $DEVICE_ID=1001
MM184 39 18 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1176 $Y=2468  $PIN_XY=1206,2470,1176,2468,1146,2470 $DEVICE_ID=1001
MM185 3 25 48 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=672 $Y=2762  $PIN_XY=702,2760,672,2762,642,2760 $DEVICE_ID=1001
MM186 3 18 40 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=672 $Y=2468  $PIN_XY=702,2470,672,2468,642,2470 $DEVICE_ID=1001
MM187 48 49 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=504 $Y=2942  $PIN_XY=534,2760,504,2942,474,2760 $DEVICE_ID=1001
MM188 40 41 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=504 $Y=2288  $PIN_XY=534,2470,504,2288,474,2470 $DEVICE_ID=1001
MM189 142 48 49 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=2942  $PIN_XY=366,2760,336,2942,306,2760 $DEVICE_ID=1001
MM190 142 40 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=2288  $PIN_XY=366,2470,336,2288,306,2470 $DEVICE_ID=1001
MM191 49 25 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=2762  $PIN_XY=198,2760,168,2762,138,2760 $DEVICE_ID=1001
MM192 41 18 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=2468  $PIN_XY=198,2470,168,2468,138,2470 $DEVICE_ID=1001
XX73A2B172155 131 130 179 188 fill_sram_inverted $T=3834 6538 1 0 $X=3810 $Y=5822
XX73A2B172156 133 132 180 189 fill_sram_inverted $T=3834 7846 1 0 $X=3810 $Y=7130
XX73A2B172157 135 134 181 190 fill_sram_inverted $T=3834 10462 1 0 $X=3810 $Y=9746
XX73A2B172158 136 137 182 191 fill_sram_inverted $T=3834 9154 1 0 $X=3810 $Y=8438
XX73A2B172159 139 138 183 192 fill_sram_inverted $T=3834 3922 1 0 $X=3810 $Y=3206
XX73A2B172160 140 141 184 193 fill_sram_inverted $T=3834 5230 1 0 $X=3810 $Y=4514
XX73A2B172161 142 143 185 194 fill_sram_inverted $T=3834 2614 1 0 $X=3810 $Y=1898
XX73A2B172162 144 145 186 195 fill_sram_inverted $T=3834 1306 1 0 $X=3810 $Y=590
XX73A2B172163 140 130 184 188 fill_sram $T=3834 5232 0 0 $X=3810 $Y=5168
XX73A2B172164 131 132 179 189 fill_sram $T=3834 6540 0 0 $X=3810 $Y=6476
XX73A2B172165 136 134 182 190 fill_sram $T=3834 9156 0 0 $X=3810 $Y=9092
XX73A2B172166 133 137 180 191 fill_sram $T=3834 7848 0 0 $X=3810 $Y=7784
XX73A2B172167 142 138 185 192 fill_sram $T=3834 2616 0 0 $X=3810 $Y=2552
XX73A2B172168 139 141 183 193 fill_sram $T=3834 3924 0 0 $X=3810 $Y=3860
XX73A2B172169 144 143 186 194 fill_sram $T=3834 1308 0 0 $X=3810 $Y=1244
XX73A2B172170 146 145 187 195 fill_sram $T=3834 0 0 0 $X=3810 $Y=-64
XX73A2B172171 2 2 3 3 4 4 5 5 6 6 7 
+	7 8 8 9 9 18 19 20 147 148 149 
+	150 151 152 153 154 34 35 36 37 38 39 
+	40 41 143 145 144 142 2 3 5 6 7 
+	4 8 9 2 3 5 6 7 4 8 9 
+	21 146 186 185 194 195 187 VCELLR4 $T=0 2614 1 0 $X=-54 $Y=-64
XX73A2B172172 2 2 3 3 4 4 5 5 6 6 7 
+	7 8 8 9 9 22 23 24 42 43 44 
+	45 46 47 48 49 50 51 52 53 54 55 
+	56 57 141 138 139 140 2 3 5 6 7 
+	4 8 9 2 3 5 6 7 4 8 9 
+	25 142 183 184 193 192 185 VCELLR4 $T=0 5230 1 0 $X=-54 $Y=2552
XX73A2B172173 2 2 3 3 4 4 5 5 6 6 7 
+	7 8 8 9 9 26 27 28 58 59 60 
+	61 62 63 64 65 66 67 68 69 70 71 
+	72 73 132 130 131 133 2 3 5 6 7 
+	4 8 9 2 3 5 6 7 4 8 9 
+	29 140 179 180 189 188 184 VCELLR4 $T=0 7846 1 0 $X=-54 $Y=5168
XX73A2B172174 2 2 3 3 4 4 5 5 6 6 7 
+	7 8 8 9 9 30 31 32 74 75 76 
+	77 78 79 80 81 163 164 165 166 167 168 
+	169 170 134 137 136 135 2 3 5 6 7 
+	4 8 9 2 3 5 6 7 4 8 9 
+	33 133 182 181 190 191 180 VCELLR4 $T=0 10462 1 0 $X=-54 $Y=7784
XX73A2B172175 10 10 11 11 12 12 13 13 14 14 15 
+	15 16 16 17 17 18 19 20 155 156 157 
+	158 159 160 161 162 82 83 84 85 86 87 
+	88 89 143 145 144 142 10 11 13 14 15 
+	12 16 17 10 11 13 14 15 12 16 17 
+	21 146 186 185 194 195 187 VCELLR4 $T=4032 2614 1 0 $X=3978 $Y=-64
XX73A2B172176 10 10 11 11 12 12 13 13 14 14 15 
+	15 16 16 17 17 22 23 24 90 91 92 
+	93 94 95 96 97 98 99 100 101 102 103 
+	104 105 141 138 139 140 10 11 13 14 15 
+	12 16 17 10 11 13 14 15 12 16 17 
+	25 142 183 184 193 192 185 VCELLR4 $T=4032 5230 1 0 $X=3978 $Y=2552
XX73A2B172177 10 10 11 11 12 12 13 13 14 14 15 
+	15 16 16 17 17 26 27 28 106 107 108 
+	109 110 111 112 113 114 115 116 117 118 119 
+	120 121 132 130 131 133 10 11 13 14 15 
+	12 16 17 10 11 13 14 15 12 16 17 
+	29 140 179 180 189 188 184 VCELLR4 $T=4032 7846 1 0 $X=3978 $Y=5168
XX73A2B172178 10 10 11 11 12 12 13 13 14 14 15 
+	15 16 16 17 17 30 31 32 122 123 124 
+	125 126 127 128 129 171 172 173 174 175 176 
+	177 178 134 137 136 135 10 11 13 14 15 
+	12 16 17 10 11 13 14 15 12 16 17 
+	33 133 182 181 190 191 180 VCELLR4 $T=4032 10462 1 0 $X=3978 $Y=7784
.ends sram_array_16r_8c

* Hierarchy Level 0

* Top of hierarchy  cell=top_level
.subckt top_level CLK A<4> WENB A<0> A<1> A<2> A<3> 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 23
+	24 D<3> Q<3> D<2> Q<2> D<1> Q<1> D<0> Q<0> 33 34
+	35 36 37 38 39 40 41 42 43 44 45
+	46 47 48 49 50 51 52 53 54 55 56
+	57 58 59 60 61 62 63 64 65 66 67
+	68 VDD! GND!
MM1 15 64 112 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11760 $Y=11624  $PIN_XY=11790,11626,11760,11624,11730,11626 $DEVICE_ID=1001
MM2 12 77 148 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11592 $Y=13313  $PIN_XY=(11622,13418,11622,13224),11592,13313,(11562,13418,11562,13224) $DEVICE_ID=1001
MM3 112 113 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11592 $Y=11444  $PIN_XY=11622,11626,11592,11444,11562,11626 $DEVICE_ID=1001
MM4 GND! 112 113 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11424 $Y=11444  $PIN_XY=11454,11626,11424,11444,11394,11626 $DEVICE_ID=1001
MM5 148 A<4> 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11256 $Y=13313  $PIN_XY=(11286,13418,11286,13224),11256,13313,(11226,13418,11226,13224) $DEVICE_ID=1001
MM6 113 64 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=11624  $PIN_XY=11286,11626,11256,11624,11226,11626 $DEVICE_ID=1001
MM7 14 64 114 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=11624  $PIN_XY=10782,11626,10752,11624,10722,11626 $DEVICE_ID=1001
MM8 15 77 149 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10584 $Y=13313  $PIN_XY=(10614,13418,10614,13224),10584,13313,(10554,13418,10554,13224) $DEVICE_ID=1001
MM9 114 115 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10584 $Y=11444  $PIN_XY=10614,11626,10584,11444,10554,11626 $DEVICE_ID=1001
MM10 GND! 114 115 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10416 $Y=11444  $PIN_XY=10446,11626,10416,11444,10386,11626 $DEVICE_ID=1001
MM11 149 A<4> 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10248 $Y=13313  $PIN_XY=(10278,13418,10278,13224),10248,13313,(10218,13418,10218,13224) $DEVICE_ID=1001
MM12 115 64 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10248 $Y=11624  $PIN_XY=10278,11626,10248,11624,10218,11626 $DEVICE_ID=1001
MM13 11 64 116 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9744 $Y=11624  $PIN_XY=9774,11626,9744,11624,9714,11626 $DEVICE_ID=1001
MM14 24 77 146 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9576 $Y=13313  $PIN_XY=(9606,13418,9606,13224),9576,13313,(9546,13418,9546,13224) $DEVICE_ID=1001
MM15 116 117 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9576 $Y=11444  $PIN_XY=9606,11626,9576,11444,9546,11626 $DEVICE_ID=1001
MM16 GND! 116 117 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9408 $Y=11444  $PIN_XY=9438,11626,9408,11444,9378,11626 $DEVICE_ID=1001
MM17 146 A<4> 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9240 $Y=13313  $PIN_XY=(9270,13418,9270,13224),9240,13313,(9210,13418,9210,13224) $DEVICE_ID=1001
MM18 117 64 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9240 $Y=11624  $PIN_XY=9270,11626,9240,11624,9210,11626 $DEVICE_ID=1001
MM19 10 64 118 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8736 $Y=11624  $PIN_XY=8766,11626,8736,11624,8706,11626 $DEVICE_ID=1001
MM20 14 77 147 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8568 $Y=13313  $PIN_XY=(8598,13418,8598,13224),8568,13313,(8538,13418,8538,13224) $DEVICE_ID=1001
MM21 118 119 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8568 $Y=11444  $PIN_XY=8598,11626,8568,11444,8538,11626 $DEVICE_ID=1001
MM22 GND! 118 119 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8400 $Y=11444  $PIN_XY=8430,11626,8400,11444,8370,11626 $DEVICE_ID=1001
MM23 147 A<4> 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8232 $Y=13313  $PIN_XY=(8262,13418,8262,13224),8232,13313,(8202,13418,8202,13224) $DEVICE_ID=1001
MM24 119 64 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=11624  $PIN_XY=8262,11626,8232,11624,8202,11626 $DEVICE_ID=1001
MM25 9 64 104 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=11624  $PIN_XY=7758,11626,7728,11624,7698,11626 $DEVICE_ID=1001
MM26 23 77 145 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7560 $Y=13313  $PIN_XY=(7590,13418,7590,13224),7560,13313,(7530,13418,7530,13224) $DEVICE_ID=1001
MM27 104 105 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7560 $Y=11444  $PIN_XY=7590,11626,7560,11444,7530,11626 $DEVICE_ID=1001
MM28 GND! 104 105 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7392 $Y=11444  $PIN_XY=7422,11626,7392,11444,7362,11626 $DEVICE_ID=1001
MM29 145 A<4> 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7224 $Y=13313  $PIN_XY=(7254,13418,7254,13224),7224,13313,(7194,13418,7194,13224) $DEVICE_ID=1001
MM30 105 64 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7224 $Y=11624  $PIN_XY=7254,11626,7224,11624,7194,11626 $DEVICE_ID=1001
MM31 13 64 106 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6720 $Y=11624  $PIN_XY=6750,11626,6720,11624,6690,11626 $DEVICE_ID=1001
MM32 11 77 144 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6552 $Y=13313  $PIN_XY=(6582,13418,6582,13224),6552,13313,(6522,13418,6522,13224) $DEVICE_ID=1001
MM33 106 107 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6552 $Y=11444  $PIN_XY=6582,11626,6552,11444,6522,11626 $DEVICE_ID=1001
MM34 GND! 106 107 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6384 $Y=11444  $PIN_XY=6414,11626,6384,11444,6354,11626 $DEVICE_ID=1001
MM35 144 A<4> 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6216 $Y=13313  $PIN_XY=(6246,13418,6246,13224),6216,13313,(6186,13418,6186,13224) $DEVICE_ID=1001
MM36 107 64 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6216 $Y=11624  $PIN_XY=6246,11626,6216,11624,6186,11626 $DEVICE_ID=1001
MM37 19 64 108 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5712 $Y=11624  $PIN_XY=5742,11626,5712,11624,5682,11626 $DEVICE_ID=1001
MM38 22 77 143 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5544 $Y=13313  $PIN_XY=(5574,13418,5574,13224),5544,13313,(5514,13418,5514,13224) $DEVICE_ID=1001
MM39 108 109 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5544 $Y=11444  $PIN_XY=5574,11626,5544,11444,5514,11626 $DEVICE_ID=1001
MM40 GND! 108 109 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5376 $Y=11444  $PIN_XY=5406,11626,5376,11444,5346,11626 $DEVICE_ID=1001
MM41 143 A<4> 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5208 $Y=13313  $PIN_XY=(5238,13418,5238,13224),5208,13313,(5178,13418,5178,13224) $DEVICE_ID=1001
MM42 109 64 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5208 $Y=11624  $PIN_XY=5238,11626,5208,11624,5178,11626 $DEVICE_ID=1001
MM43 17 64 110 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4704 $Y=11624  $PIN_XY=4734,11626,4704,11624,4674,11626 $DEVICE_ID=1001
MM44 10 77 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4536 $Y=13313  $PIN_XY=(4566,13418,4566,13224),4536,13313,(4506,13418,4506,13224) $DEVICE_ID=1001
MM45 110 111 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4536 $Y=11444  $PIN_XY=4566,11626,4536,11444,4506,11626 $DEVICE_ID=1001
MM46 GND! 110 111 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4368 $Y=11444  $PIN_XY=4398,11626,4368,11444,4338,11626 $DEVICE_ID=1001
MM47 142 A<4> 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4200 $Y=13313  $PIN_XY=(4230,13418,4230,13224),4200,13313,(4170,13418,4170,13224) $DEVICE_ID=1001
MM48 111 64 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=11624  $PIN_XY=4230,11626,4200,11624,4170,11626 $DEVICE_ID=1001
MM49 GND! 85 64 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=11444  $PIN_XY=3894,11626,3864,11444,3834,11626 $DEVICE_ID=1001
MM50 GND! 76 63 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=10790  $PIN_XY=3894,10608,3864,10790,3834,10608 $DEVICE_ID=1001
MM51 GND! 84 62 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=10136  $PIN_XY=3894,10318,3864,10136,3834,10318 $DEVICE_ID=1001
MM52 GND! 75 61 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=9482  $PIN_XY=3894,9300,3864,9482,3834,9300 $DEVICE_ID=1001
MM53 GND! 83 60 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=8828  $PIN_XY=3894,9010,3864,8828,3834,9010 $DEVICE_ID=1001
MM54 GND! 74 59 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=8174  $PIN_XY=3894,7992,3864,8174,3834,7992 $DEVICE_ID=1001
MM55 GND! 78 58 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=7520  $PIN_XY=3894,7702,3864,7520,3834,7702 $DEVICE_ID=1001
MM56 GND! 69 57 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=6866  $PIN_XY=3894,6684,3864,6866,3834,6684 $DEVICE_ID=1001
MM57 GND! 79 56 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=6212  $PIN_XY=3894,6394,3864,6212,3834,6394 $DEVICE_ID=1001
MM58 GND! 70 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=5558  $PIN_XY=3894,5376,3864,5558,3834,5376 $DEVICE_ID=1001
MM59 GND! 80 54 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=4904  $PIN_XY=3894,5086,3864,4904,3834,5086 $DEVICE_ID=1001
MM60 GND! 71 53 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=4250  $PIN_XY=3894,4068,3864,4250,3834,4068 $DEVICE_ID=1001
MM61 64 85 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=11444  $PIN_XY=3726,11626,3696,11444,3666,11626 $DEVICE_ID=1001
MM62 63 76 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=10790  $PIN_XY=3726,10608,3696,10790,3666,10608 $DEVICE_ID=1001
MM63 62 84 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=10136  $PIN_XY=3726,10318,3696,10136,3666,10318 $DEVICE_ID=1001
MM64 61 75 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=9482  $PIN_XY=3726,9300,3696,9482,3666,9300 $DEVICE_ID=1001
MM65 60 83 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=8828  $PIN_XY=3726,9010,3696,8828,3666,9010 $DEVICE_ID=1001
MM66 59 74 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=8174  $PIN_XY=3726,7992,3696,8174,3666,7992 $DEVICE_ID=1001
MM67 58 78 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=7520  $PIN_XY=3726,7702,3696,7520,3666,7702 $DEVICE_ID=1001
MM68 57 69 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=6866  $PIN_XY=3726,6684,3696,6866,3666,6684 $DEVICE_ID=1001
MM69 56 79 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=6212  $PIN_XY=3726,6394,3696,6212,3666,6394 $DEVICE_ID=1001
MM70 55 70 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=5558  $PIN_XY=3726,5376,3696,5558,3666,5376 $DEVICE_ID=1001
MM71 54 80 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=4904  $PIN_XY=3726,5086,3696,4904,3666,5086 $DEVICE_ID=1001
MM72 53 71 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=4250  $PIN_XY=3726,4068,3696,4250,3666,4068 $DEVICE_ID=1001
MM73 GND! 46 85 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=11444  $PIN_XY=3390,11626,3360,11444,3330,11626 $DEVICE_ID=1001
MM74 GND! 48 76 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=10790  $PIN_XY=3390,10608,3360,10790,3330,10608 $DEVICE_ID=1001
MM75 GND! 45 84 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=10136  $PIN_XY=3390,10318,3360,10136,3330,10318 $DEVICE_ID=1001
MM76 GND! 47 75 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=9482  $PIN_XY=3390,9300,3360,9482,3330,9300 $DEVICE_ID=1001
MM77 GND! 41 83 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=8828  $PIN_XY=3390,9010,3360,8828,3330,9010 $DEVICE_ID=1001
MM78 GND! 44 74 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=8174  $PIN_XY=3390,7992,3360,8174,3330,7992 $DEVICE_ID=1001
MM79 GND! 40 78 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=7520  $PIN_XY=3390,7702,3360,7520,3330,7702 $DEVICE_ID=1001
MM80 GND! 43 69 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=6866  $PIN_XY=3390,6684,3360,6866,3330,6684 $DEVICE_ID=1001
MM81 GND! 39 79 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=6212  $PIN_XY=3390,6394,3360,6212,3330,6394 $DEVICE_ID=1001
MM82 GND! 42 70 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=5558  $PIN_XY=3390,5376,3360,5558,3330,5376 $DEVICE_ID=1001
MM83 GND! 35 80 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=4904  $PIN_XY=3390,5086,3360,4904,3330,5086 $DEVICE_ID=1001
MM84 GND! 38 71 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=4250  $PIN_XY=3390,4068,3360,4250,3330,4068 $DEVICE_ID=1001
MM85 85 46 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=11444  $PIN_XY=3222,11626,3192,11444,3162,11626 $DEVICE_ID=1001
MM86 76 48 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=10790  $PIN_XY=3222,10608,3192,10790,3162,10608 $DEVICE_ID=1001
MM87 84 45 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=10136  $PIN_XY=3222,10318,3192,10136,3162,10318 $DEVICE_ID=1001
MM88 75 47 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=9482  $PIN_XY=3222,9300,3192,9482,3162,9300 $DEVICE_ID=1001
MM89 83 41 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=8828  $PIN_XY=3222,9010,3192,8828,3162,9010 $DEVICE_ID=1001
MM90 74 44 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=8174  $PIN_XY=3222,7992,3192,8174,3162,7992 $DEVICE_ID=1001
MM91 78 40 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=7520  $PIN_XY=3222,7702,3192,7520,3162,7702 $DEVICE_ID=1001
MM92 69 43 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=6866  $PIN_XY=3222,6684,3192,6866,3162,6684 $DEVICE_ID=1001
MM93 79 39 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=6212  $PIN_XY=3222,6394,3192,6212,3162,6394 $DEVICE_ID=1001
MM94 70 42 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=5558  $PIN_XY=3222,5376,3192,5558,3162,5376 $DEVICE_ID=1001
MM95 80 35 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=4904  $PIN_XY=3222,5086,3192,4904,3162,5086 $DEVICE_ID=1001
MM96 71 38 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=4250  $PIN_XY=3222,4068,3192,4250,3162,4068 $DEVICE_ID=1001
MM97 15 49 96 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11760 $Y=1454  $PIN_XY=11790,1452,11760,1454,11730,1452 $DEVICE_ID=1001
MM98 96 97 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11592 $Y=1634  $PIN_XY=11622,1452,11592,1634,11562,1452 $DEVICE_ID=1001
MM99 GND! 96 97 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11424 $Y=1634  $PIN_XY=11454,1452,11424,1634,11394,1452 $DEVICE_ID=1001
MM100 97 49 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=1454  $PIN_XY=11286,1452,11256,1454,11226,1452 $DEVICE_ID=1001
MM101 15 WENB 151 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11256 $Y=1073  $PIN_XY=11286,1162,11256,1073,11226,1162 $DEVICE_ID=1001
MM102 151 87 68 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11088 $Y=1073  $PIN_XY=11118,1162,11088,1073,11058,1162 $DEVICE_ID=1001
MM103 68 A<4> 150 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10920 $Y=1073  $PIN_XY=10950,1162,10920,1073,10890,1162 $DEVICE_ID=1001
MM104 14 49 98 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=1454  $PIN_XY=10782,1452,10752,1454,10722,1452 $DEVICE_ID=1001
MM105 150 WENB 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10752 $Y=1073  $PIN_XY=10782,1162,10752,1073,10722,1162 $DEVICE_ID=1001
MM106 98 99 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10584 $Y=1634  $PIN_XY=10614,1452,10584,1634,10554,1452 $DEVICE_ID=1001
MM107 GND! 98 99 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10416 $Y=1634  $PIN_XY=10446,1452,10416,1634,10386,1452 $DEVICE_ID=1001
MM108 99 49 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10248 $Y=1454  $PIN_XY=10278,1452,10248,1454,10218,1452 $DEVICE_ID=1001
MM109 11 49 100 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9744 $Y=1454  $PIN_XY=9774,1452,9744,1454,9714,1452 $DEVICE_ID=1001
MM110 100 101 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9576 $Y=1634  $PIN_XY=9606,1452,9576,1634,9546,1452 $DEVICE_ID=1001
MM111 GND! 100 101 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9408 $Y=1634  $PIN_XY=9438,1452,9408,1634,9378,1452 $DEVICE_ID=1001
MM112 101 49 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9240 $Y=1454  $PIN_XY=9270,1452,9240,1454,9210,1452 $DEVICE_ID=1001
MM113 14 WENB 153 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9240 $Y=1073  $PIN_XY=9270,1162,9240,1073,9210,1162 $DEVICE_ID=1001
MM114 153 87 67 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9072 $Y=1073  $PIN_XY=9102,1162,9072,1073,9042,1162 $DEVICE_ID=1001
MM115 67 A<4> 152 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8904 $Y=1073  $PIN_XY=8934,1162,8904,1073,8874,1162 $DEVICE_ID=1001
MM116 10 49 102 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8736 $Y=1454  $PIN_XY=8766,1452,8736,1454,8706,1452 $DEVICE_ID=1001
MM117 152 WENB 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8736 $Y=1073  $PIN_XY=8766,1162,8736,1073,8706,1162 $DEVICE_ID=1001
MM118 102 103 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8568 $Y=1634  $PIN_XY=8598,1452,8568,1634,8538,1452 $DEVICE_ID=1001
MM119 GND! 102 103 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8400 $Y=1634  $PIN_XY=8430,1452,8400,1634,8370,1452 $DEVICE_ID=1001
MM120 103 49 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=1454  $PIN_XY=8262,1452,8232,1454,8202,1452 $DEVICE_ID=1001
MM121 9 49 88 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=1454  $PIN_XY=7758,1452,7728,1454,7698,1452 $DEVICE_ID=1001
MM122 88 89 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7560 $Y=1634  $PIN_XY=7590,1452,7560,1634,7530,1452 $DEVICE_ID=1001
MM123 GND! 88 89 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7392 $Y=1634  $PIN_XY=7422,1452,7392,1634,7362,1452 $DEVICE_ID=1001
MM124 89 49 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7224 $Y=1454  $PIN_XY=7254,1452,7224,1454,7194,1452 $DEVICE_ID=1001
MM125 11 WENB 155 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7224 $Y=1073  $PIN_XY=7254,1162,7224,1073,7194,1162 $DEVICE_ID=1001
MM126 155 87 66 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7056 $Y=1073  $PIN_XY=7086,1162,7056,1073,7026,1162 $DEVICE_ID=1001
MM127 66 A<4> 154 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6888 $Y=1073  $PIN_XY=6918,1162,6888,1073,6858,1162 $DEVICE_ID=1001
MM128 13 49 90 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6720 $Y=1454  $PIN_XY=6750,1452,6720,1454,6690,1452 $DEVICE_ID=1001
MM129 154 WENB 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6720 $Y=1073  $PIN_XY=6750,1162,6720,1073,6690,1162 $DEVICE_ID=1001
MM130 90 91 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6552 $Y=1634  $PIN_XY=6582,1452,6552,1634,6522,1452 $DEVICE_ID=1001
MM131 GND! 90 91 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6384 $Y=1634  $PIN_XY=6414,1452,6384,1634,6354,1452 $DEVICE_ID=1001
MM132 91 49 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6216 $Y=1454  $PIN_XY=6246,1452,6216,1454,6186,1452 $DEVICE_ID=1001
MM133 19 49 92 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5712 $Y=1454  $PIN_XY=5742,1452,5712,1454,5682,1452 $DEVICE_ID=1001
MM134 92 93 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5544 $Y=1634  $PIN_XY=5574,1452,5544,1634,5514,1452 $DEVICE_ID=1001
MM135 GND! 92 93 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5376 $Y=1634  $PIN_XY=5406,1452,5376,1634,5346,1452 $DEVICE_ID=1001
MM136 10 WENB 157 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5376 $Y=1073  $PIN_XY=5406,1162,5376,1073,5346,1162 $DEVICE_ID=1001
MM137 93 49 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5208 $Y=1454  $PIN_XY=5238,1452,5208,1454,5178,1452 $DEVICE_ID=1001
MM138 157 87 65 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5208 $Y=1073  $PIN_XY=5238,1162,5208,1073,5178,1162 $DEVICE_ID=1001
MM139 65 A<4> 156 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5040 $Y=1073  $PIN_XY=5070,1162,5040,1073,5010,1162 $DEVICE_ID=1001
MM140 156 WENB 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4872 $Y=1073  $PIN_XY=4902,1162,4872,1073,4842,1162 $DEVICE_ID=1001
MM141 17 49 94 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4704 $Y=1454  $PIN_XY=4734,1452,4704,1454,4674,1452 $DEVICE_ID=1001
MM142 94 95 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4536 $Y=1634  $PIN_XY=4566,1452,4536,1634,4506,1452 $DEVICE_ID=1001
MM143 GND! 94 95 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4368 $Y=1634  $PIN_XY=4398,1452,4368,1634,4338,1452 $DEVICE_ID=1001
MM144 95 49 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=1454  $PIN_XY=4230,1452,4200,1454,4170,1452 $DEVICE_ID=1001
MM145 GND! 81 52 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=3596  $PIN_XY=3894,3778,3864,3596,3834,3778 $DEVICE_ID=1001
MM146 GND! 72 51 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=2942  $PIN_XY=3894,2760,3864,2942,3834,2760 $DEVICE_ID=1001
MM147 GND! 82 50 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=2288  $PIN_XY=3894,2470,3864,2288,3834,2470 $DEVICE_ID=1001
MM148 GND! 73 49 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=1634  $PIN_XY=3894,1452,3864,1634,3834,1452 $DEVICE_ID=1001
MM149 GND! A<4> 87 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=980  $PIN_XY=3894,1162,3864,980,3834,1162 $DEVICE_ID=1001
MM150 52 81 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=3596  $PIN_XY=3726,3778,3696,3596,3666,3778 $DEVICE_ID=1001
MM151 51 72 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=2942  $PIN_XY=3726,2760,3696,2942,3666,2760 $DEVICE_ID=1001
MM152 50 82 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=2288  $PIN_XY=3726,2470,3696,2288,3666,2470 $DEVICE_ID=1001
MM153 49 73 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=1634  $PIN_XY=3726,1452,3696,1634,3666,1452 $DEVICE_ID=1001
MM154 87 A<4> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=980  $PIN_XY=3726,1162,3696,980,3666,1162 $DEVICE_ID=1001
MM155 GND! 34 81 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=3596  $PIN_XY=3390,3778,3360,3596,3330,3778 $DEVICE_ID=1001
MM156 GND! 37 72 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=2942  $PIN_XY=3390,2760,3360,2942,3330,2760 $DEVICE_ID=1001
MM157 GND! 33 82 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=2288  $PIN_XY=3390,2470,3360,2288,3330,2470 $DEVICE_ID=1001
MM158 GND! 36 73 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=1634  $PIN_XY=3390,1452,3360,1634,3330,1452 $DEVICE_ID=1001
MM159 81 34 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=3596  $PIN_XY=3222,3778,3192,3596,3162,3778 $DEVICE_ID=1001
MM160 72 37 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=2942  $PIN_XY=3222,2760,3192,2942,3162,2760 $DEVICE_ID=1001
MM161 82 33 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=2288  $PIN_XY=3222,2470,3192,2288,3162,2470 $DEVICE_ID=1001
MM162 73 36 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=1634  $PIN_XY=3222,1452,3192,1634,3162,1452 $DEVICE_ID=1001
MM163 36 A<3> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2856 $Y=1454  $PIN_XY=2886,1452,2856,1454,2826,1452 $DEVICE_ID=1001
MM164 36 A<2> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2520 $Y=1454  $PIN_XY=2550,1452,2520,1454,2490,1452 $DEVICE_ID=1001
MM165 36 A<1> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2184 $Y=1454  $PIN_XY=2214,1452,2184,1454,2154,1452 $DEVICE_ID=1001
MM166 36 A<0> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1848 $Y=1454  $PIN_XY=1878,1452,1848,1454,1818,1452 $DEVICE_ID=1001
MM167 33 A<3> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1512 $Y=1454  $PIN_XY=1542,1452,1512,1454,1482,1452 $DEVICE_ID=1001
MM168 33 A<2> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1176 $Y=1454  $PIN_XY=1206,1452,1176,1454,1146,1452 $DEVICE_ID=1001
MM169 33 A<1> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=840 $Y=1454  $PIN_XY=870,1452,840,1454,810,1452 $DEVICE_ID=1001
MM170 33 86 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=504 $Y=1454  $PIN_XY=534,1452,504,1454,474,1452 $DEVICE_ID=1001
MM171 VDD! 120 Q<0> pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=11424 $Y=326  $PIN_XY=(11454,508,11454,338),11424,326,(11394,508,11394,338) $DEVICE_ID=1003
MM172 Q<0> 120 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=11256 $Y=326  $PIN_XY=(11286,508,11286,338),11256,326,(11226,508,11226,338) $DEVICE_ID=1003
MM173 VDD! 68 120 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=10920 $Y=326  $PIN_XY=(10950,508,10950,338),10920,326,(10890,508,10890,338) $DEVICE_ID=1003
MM174 120 68 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=10752 $Y=326  $PIN_XY=(10782,508,10782,338),10752,326,(10722,508,10722,338) $DEVICE_ID=1003
MM175 VDD! 121 Q<1> pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=9408 $Y=326  $PIN_XY=(9438,508,9438,338),9408,326,(9378,508,9378,338) $DEVICE_ID=1003
MM176 Q<1> 121 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=9240 $Y=326  $PIN_XY=(9270,508,9270,338),9240,326,(9210,508,9210,338) $DEVICE_ID=1003
MM177 VDD! 67 121 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=8904 $Y=326  $PIN_XY=(8934,508,8934,338),8904,326,(8874,508,8874,338) $DEVICE_ID=1003
MM178 121 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=8736 $Y=326  $PIN_XY=(8766,508,8766,338),8736,326,(8706,508,8706,338) $DEVICE_ID=1003
MM179 VDD! 122 Q<2> pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=7392 $Y=326  $PIN_XY=(7422,508,7422,338),7392,326,(7362,508,7362,338) $DEVICE_ID=1003
MM180 Q<2> 122 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=7224 $Y=326  $PIN_XY=(7254,508,7254,338),7224,326,(7194,508,7194,338) $DEVICE_ID=1003
MM181 VDD! 66 122 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=6888 $Y=326  $PIN_XY=(6918,508,6918,338),6888,326,(6858,508,6858,338) $DEVICE_ID=1003
MM182 122 66 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=6720 $Y=326  $PIN_XY=(6750,508,6750,338),6720,326,(6690,508,6690,338) $DEVICE_ID=1003
MM183 VDD! 123 Q<3> pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=5544 $Y=326  $PIN_XY=(5574,508,5574,338),5544,326,(5514,508,5514,338) $DEVICE_ID=1003
MM184 Q<3> 123 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=5376 $Y=326  $PIN_XY=(5406,508,5406,338),5376,326,(5346,508,5346,338) $DEVICE_ID=1003
MM185 VDD! 65 123 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=5040 $Y=326  $PIN_XY=(5070,508,5070,338),5040,326,(5010,508,5010,338) $DEVICE_ID=1003
MM186 123 65 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=4872 $Y=326  $PIN_XY=(4902,508,4902,338),4872,326,(4842,508,4842,338) $DEVICE_ID=1003
MM187 VDD! 85 64 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=11444  $PIN_XY=(3894,11432,3894,11262),3864,11444,(3834,11432,3834,11262) $DEVICE_ID=1003
MM188 VDD! 76 63 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=10790  $PIN_XY=(3894,10972,3894,10802),3864,10790,(3834,10972,3834,10802) $DEVICE_ID=1003
MM189 VDD! 84 62 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=10136  $PIN_XY=(3894,10124,3894,9954),3864,10136,(3834,10124,3834,9954) $DEVICE_ID=1003
MM190 VDD! 75 61 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=9482  $PIN_XY=(3894,9664,3894,9494),3864,9482,(3834,9664,3834,9494) $DEVICE_ID=1003
MM191 VDD! 83 60 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=8828  $PIN_XY=(3894,8816,3894,8646),3864,8828,(3834,8816,3834,8646) $DEVICE_ID=1003
MM192 VDD! 74 59 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=8174  $PIN_XY=(3894,8356,3894,8186),3864,8174,(3834,8356,3834,8186) $DEVICE_ID=1003
MM193 VDD! 78 58 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=7520  $PIN_XY=(3894,7508,3894,7338),3864,7520,(3834,7508,3834,7338) $DEVICE_ID=1003
MM194 VDD! 69 57 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=6866  $PIN_XY=(3894,7048,3894,6878),3864,6866,(3834,7048,3834,6878) $DEVICE_ID=1003
MM195 VDD! 79 56 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=6212  $PIN_XY=(3894,6200,3894,6030),3864,6212,(3834,6200,3834,6030) $DEVICE_ID=1003
MM196 VDD! 70 55 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=5558  $PIN_XY=(3894,5740,3894,5570),3864,5558,(3834,5740,3834,5570) $DEVICE_ID=1003
MM197 VDD! 80 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=4904  $PIN_XY=(3894,4892,3894,4722),3864,4904,(3834,4892,3834,4722) $DEVICE_ID=1003
MM198 VDD! 71 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=4250  $PIN_XY=(3894,4432,3894,4262),3864,4250,(3834,4432,3834,4262) $DEVICE_ID=1003
MM199 VDD! 81 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=3596  $PIN_XY=(3894,3584,3894,3414),3864,3596,(3834,3584,3834,3414) $DEVICE_ID=1003
MM200 VDD! 72 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=2942  $PIN_XY=(3894,3124,3894,2954),3864,2942,(3834,3124,3834,2954) $DEVICE_ID=1003
MM201 VDD! 82 50 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=2288  $PIN_XY=(3894,2276,3894,2106),3864,2288,(3834,2276,3834,2106) $DEVICE_ID=1003
MM202 VDD! 73 49 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3864 $Y=1634  $PIN_XY=(3894,1816,3894,1646),3864,1634,(3834,1816,3834,1646) $DEVICE_ID=1003
MM203 VDD! A<4> 87 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3864 $Y=980  $PIN_XY=3894,798,3864,980,3834,798 $DEVICE_ID=1003
MM204 64 85 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=11444  $PIN_XY=(3726,11432,3726,11262),3696,11444,(3666,11432,3666,11262) $DEVICE_ID=1003
MM205 63 76 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=10790  $PIN_XY=(3726,10972,3726,10802),3696,10790,(3666,10972,3666,10802) $DEVICE_ID=1003
MM206 62 84 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=10136  $PIN_XY=(3726,10124,3726,9954),3696,10136,(3666,10124,3666,9954) $DEVICE_ID=1003
MM207 61 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=9482  $PIN_XY=(3726,9664,3726,9494),3696,9482,(3666,9664,3666,9494) $DEVICE_ID=1003
MM208 60 83 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=8828  $PIN_XY=(3726,8816,3726,8646),3696,8828,(3666,8816,3666,8646) $DEVICE_ID=1003
MM209 59 74 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=8174  $PIN_XY=(3726,8356,3726,8186),3696,8174,(3666,8356,3666,8186) $DEVICE_ID=1003
MM210 58 78 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=7520  $PIN_XY=(3726,7508,3726,7338),3696,7520,(3666,7508,3666,7338) $DEVICE_ID=1003
MM211 57 69 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=6866  $PIN_XY=(3726,7048,3726,6878),3696,6866,(3666,7048,3666,6878) $DEVICE_ID=1003
MM212 56 79 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=6212  $PIN_XY=(3726,6200,3726,6030),3696,6212,(3666,6200,3666,6030) $DEVICE_ID=1003
MM213 55 70 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=5558  $PIN_XY=(3726,5740,3726,5570),3696,5558,(3666,5740,3666,5570) $DEVICE_ID=1003
MM214 54 80 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=4904  $PIN_XY=(3726,4892,3726,4722),3696,4904,(3666,4892,3666,4722) $DEVICE_ID=1003
MM215 53 71 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=4250  $PIN_XY=(3726,4432,3726,4262),3696,4250,(3666,4432,3666,4262) $DEVICE_ID=1003
MM216 52 81 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=3596  $PIN_XY=(3726,3584,3726,3414),3696,3596,(3666,3584,3666,3414) $DEVICE_ID=1003
MM217 51 72 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=2942  $PIN_XY=(3726,3124,3726,2954),3696,2942,(3666,3124,3666,2954) $DEVICE_ID=1003
MM218 50 82 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=2288  $PIN_XY=(3726,2276,3726,2106),3696,2288,(3666,2276,3666,2106) $DEVICE_ID=1003
MM219 49 73 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3696 $Y=1634  $PIN_XY=(3726,1816,3726,1646),3696,1634,(3666,1816,3666,1646) $DEVICE_ID=1003
MM220 87 A<4> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3696 $Y=980  $PIN_XY=3726,798,3696,980,3666,798 $DEVICE_ID=1003
MM221 VDD! 46 85 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=11444  $PIN_XY=(3390,11432,3390,11262),3360,11444,(3330,11432,3330,11262) $DEVICE_ID=1003
MM222 VDD! 48 76 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=10790  $PIN_XY=(3390,10972,3390,10802),3360,10790,(3330,10972,3330,10802) $DEVICE_ID=1003
MM223 VDD! 45 84 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=10136  $PIN_XY=(3390,10124,3390,9954),3360,10136,(3330,10124,3330,9954) $DEVICE_ID=1003
MM224 VDD! 47 75 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=9482  $PIN_XY=(3390,9664,3390,9494),3360,9482,(3330,9664,3330,9494) $DEVICE_ID=1003
MM225 VDD! 41 83 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=8828  $PIN_XY=(3390,8816,3390,8646),3360,8828,(3330,8816,3330,8646) $DEVICE_ID=1003
MM226 VDD! 44 74 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=8174  $PIN_XY=(3390,8356,3390,8186),3360,8174,(3330,8356,3330,8186) $DEVICE_ID=1003
MM227 VDD! 40 78 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=7520  $PIN_XY=(3390,7508,3390,7338),3360,7520,(3330,7508,3330,7338) $DEVICE_ID=1003
MM228 VDD! 43 69 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=6866  $PIN_XY=(3390,7048,3390,6878),3360,6866,(3330,7048,3330,6878) $DEVICE_ID=1003
MM229 VDD! 39 79 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=6212  $PIN_XY=(3390,6200,3390,6030),3360,6212,(3330,6200,3330,6030) $DEVICE_ID=1003
MM230 VDD! 42 70 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=5558  $PIN_XY=(3390,5740,3390,5570),3360,5558,(3330,5740,3330,5570) $DEVICE_ID=1003
MM231 VDD! 35 80 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=4904  $PIN_XY=(3390,4892,3390,4722),3360,4904,(3330,4892,3330,4722) $DEVICE_ID=1003
MM232 VDD! 38 71 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=4250  $PIN_XY=(3390,4432,3390,4262),3360,4250,(3330,4432,3330,4262) $DEVICE_ID=1003
MM233 VDD! 34 81 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=3596  $PIN_XY=(3390,3584,3390,3414),3360,3596,(3330,3584,3330,3414) $DEVICE_ID=1003
MM234 VDD! 37 72 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=2942  $PIN_XY=(3390,3124,3390,2954),3360,2942,(3330,3124,3330,2954) $DEVICE_ID=1003
MM235 VDD! 33 82 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=2288  $PIN_XY=(3390,2276,3390,2106),3360,2288,(3330,2276,3330,2106) $DEVICE_ID=1003
MM236 VDD! 36 73 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3360 $Y=1634  $PIN_XY=(3390,1816,3390,1646),3360,1634,(3330,1816,3330,1646) $DEVICE_ID=1003
MM237 85 46 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=11444  $PIN_XY=(3222,11432,3222,11262),3192,11444,(3162,11432,3162,11262) $DEVICE_ID=1003
MM238 76 48 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=10790  $PIN_XY=(3222,10972,3222,10802),3192,10790,(3162,10972,3162,10802) $DEVICE_ID=1003
MM239 84 45 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=10136  $PIN_XY=(3222,10124,3222,9954),3192,10136,(3162,10124,3162,9954) $DEVICE_ID=1003
MM240 75 47 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=9482  $PIN_XY=(3222,9664,3222,9494),3192,9482,(3162,9664,3162,9494) $DEVICE_ID=1003
MM241 83 41 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=8828  $PIN_XY=(3222,8816,3222,8646),3192,8828,(3162,8816,3162,8646) $DEVICE_ID=1003
MM242 74 44 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=8174  $PIN_XY=(3222,8356,3222,8186),3192,8174,(3162,8356,3162,8186) $DEVICE_ID=1003
MM243 78 40 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=7520  $PIN_XY=(3222,7508,3222,7338),3192,7520,(3162,7508,3162,7338) $DEVICE_ID=1003
MM244 69 43 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=6866  $PIN_XY=(3222,7048,3222,6878),3192,6866,(3162,7048,3162,6878) $DEVICE_ID=1003
MM245 79 39 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=6212  $PIN_XY=(3222,6200,3222,6030),3192,6212,(3162,6200,3162,6030) $DEVICE_ID=1003
MM246 70 42 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=5558  $PIN_XY=(3222,5740,3222,5570),3192,5558,(3162,5740,3162,5570) $DEVICE_ID=1003
MM247 80 35 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=4904  $PIN_XY=(3222,4892,3222,4722),3192,4904,(3162,4892,3162,4722) $DEVICE_ID=1003
MM248 71 38 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=4250  $PIN_XY=(3222,4432,3222,4262),3192,4250,(3162,4432,3162,4262) $DEVICE_ID=1003
MM249 81 34 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=3596  $PIN_XY=(3222,3584,3222,3414),3192,3596,(3162,3584,3162,3414) $DEVICE_ID=1003
MM250 72 37 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=2942  $PIN_XY=(3222,3124,3222,2954),3192,2942,(3162,3124,3162,2954) $DEVICE_ID=1003
MM251 82 33 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=2288  $PIN_XY=(3222,2276,3222,2106),3192,2288,(3162,2276,3162,2106) $DEVICE_ID=1003
MM252 73 36 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3192 $Y=1634  $PIN_XY=(3222,1816,3222,1646),3192,1634,(3162,1816,3162,1646) $DEVICE_ID=1003
MM253 VDD! A<3> 140 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=2856 $Y=12098  $PIN_XY=(2886,12280,2886,12110),2856,12098,(2826,12280,2826,12110) $DEVICE_ID=1003
MM254 140 A<3> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=2688 $Y=12098  $PIN_XY=(2718,12280,2718,12110),2688,12098,(2658,12280,2658,12110) $DEVICE_ID=1003
MM255 VDD! A<2> 141 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=2184 $Y=12098  $PIN_XY=(2214,12280,2214,12110),2184,12098,(2154,12280,2154,12110) $DEVICE_ID=1003
MM256 141 A<2> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=2016 $Y=12098  $PIN_XY=(2046,12280,2046,12110),2016,12098,(1986,12280,1986,12110) $DEVICE_ID=1003
MM257 VDD! A<1> 139 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=1344 $Y=12098  $PIN_XY=(1374,12280,1374,12110),1344,12098,(1314,12280,1314,12110) $DEVICE_ID=1003
MM258 139 A<1> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=1176 $Y=12098  $PIN_XY=(1206,12280,1206,12110),1176,12098,(1146,12280,1146,12110) $DEVICE_ID=1003
MM259 VDD! A<0> 86 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=672 $Y=12098  $PIN_XY=(702,12280,702,12110),672,12098,(642,12280,642,12110) $DEVICE_ID=1003
MM260 86 A<0> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=504 $Y=12098  $PIN_XY=(534,12280,534,12110),504,12098,(474,12280,474,12110) $DEVICE_ID=1003
XX73A2B1721_1 GND! VDD! 126 158 fill_sram_column_decoder_write $T=306 13080 0 0 $X=282 $Y=13016
XX73A2B1721_2 GND! VDD! 126 158 fill_sram_column_decoder_write $T=474 13080 0 0 $X=450 $Y=13016
XX73A2B1721_3 GND! VDD! 126 158 fill_sram_column_decoder_write $T=642 13080 0 0 $X=618 $Y=13016
XX73A2B1721_4 GND! VDD! 126 158 fill_sram_column_decoder_write $T=810 13080 0 0 $X=786 $Y=13016
XX73A2B1721_5 GND! VDD! 126 158 fill_sram_column_decoder_write $T=978 13080 0 0 $X=954 $Y=13016
XX73A2B1721_6 GND! VDD! 126 158 fill_sram_column_decoder_write $T=1146 13080 0 0 $X=1122 $Y=13016
XX73A2B1721_7 GND! VDD! 126 158 fill_sram_column_decoder_write $T=1314 13080 0 0 $X=1290 $Y=13016
XX73A2B1721_8 GND! VDD! 126 158 fill_sram_column_decoder_write $T=1482 13080 0 0 $X=1458 $Y=13016
XX73A2B1721_9 GND! VDD! 126 158 fill_sram_column_decoder_write $T=1650 13080 0 0 $X=1626 $Y=13016
XX73A2B1721_10 GND! VDD! 126 158 fill_sram_column_decoder_write $T=1818 13080 0 0 $X=1794 $Y=13016
XX73A2B1721_11 GND! VDD! 126 158 fill_sram_column_decoder_write $T=1986 13080 0 0 $X=1962 $Y=13016
XX73A2B1721_12 GND! VDD! 126 158 fill_sram_column_decoder_write $T=2154 13080 0 0 $X=2130 $Y=13016
XX73A2B1721_13 GND! VDD! 126 158 fill_sram_column_decoder_write $T=2322 13080 0 0 $X=2298 $Y=13016
XX73A2B1721_14 GND! VDD! 126 158 fill_sram_column_decoder_write $T=2490 13080 0 0 $X=2466 $Y=13016
XX73A2B1721_15 GND! VDD! 126 158 fill_sram_column_decoder_write $T=2658 13080 0 0 $X=2634 $Y=13016
XX73A2B1721_16 GND! VDD! 126 158 fill_sram_column_decoder_write $T=2826 13080 0 0 $X=2802 $Y=13016
XX73A2B1721_17 GND! VDD! 126 158 fill_sram_column_decoder_write $T=2994 13080 0 0 $X=2970 $Y=13016
XX73A2B1721_18 GND! VDD! 126 158 fill_sram_column_decoder_write $T=3162 13080 0 0 $X=3138 $Y=13016
XX73A2B1721_19 GND! VDD! 126 158 fill_sram_column_decoder_write $T=3330 13080 0 0 $X=3306 $Y=13016
XX73A2B17220_1 GND! VDD! 127 159 fill_sram_inverted $T=306 1306 1 0 $X=282 $Y=590
XX73A2B17220_2 GND! VDD! 127 159 fill_sram_inverted $T=474 1306 1 0 $X=450 $Y=590
XX73A2B17220_3 GND! VDD! 127 159 fill_sram_inverted $T=642 1306 1 0 $X=618 $Y=590
XX73A2B17220_4 GND! VDD! 127 159 fill_sram_inverted $T=810 1306 1 0 $X=786 $Y=590
XX73A2B17220_5 GND! VDD! 127 159 fill_sram_inverted $T=978 1306 1 0 $X=954 $Y=590
XX73A2B17220_6 GND! VDD! 127 159 fill_sram_inverted $T=1146 1306 1 0 $X=1122 $Y=590
XX73A2B17220_7 GND! VDD! 127 159 fill_sram_inverted $T=1314 1306 1 0 $X=1290 $Y=590
XX73A2B17220_8 GND! VDD! 127 159 fill_sram_inverted $T=1482 1306 1 0 $X=1458 $Y=590
XX73A2B17220_9 GND! VDD! 127 159 fill_sram_inverted $T=1650 1306 1 0 $X=1626 $Y=590
XX73A2B17220_10 GND! VDD! 127 159 fill_sram_inverted $T=1818 1306 1 0 $X=1794 $Y=590
XX73A2B17220_11 GND! VDD! 127 159 fill_sram_inverted $T=1986 1306 1 0 $X=1962 $Y=590
XX73A2B17220_12 GND! VDD! 127 159 fill_sram_inverted $T=2154 1306 1 0 $X=2130 $Y=590
XX73A2B17220_13 GND! VDD! 127 159 fill_sram_inverted $T=2322 1306 1 0 $X=2298 $Y=590
XX73A2B17220_14 GND! VDD! 127 159 fill_sram_inverted $T=2490 1306 1 0 $X=2466 $Y=590
XX73A2B17220_15 GND! VDD! 127 159 fill_sram_inverted $T=2658 1306 1 0 $X=2634 $Y=590
XX73A2B17220_16 GND! VDD! 127 159 fill_sram_inverted $T=2826 1306 1 0 $X=2802 $Y=590
XX73A2B17220_17 GND! VDD! 127 159 fill_sram_inverted $T=2994 1306 1 0 $X=2970 $Y=590
XX73A2B17220_18 GND! VDD! 127 159 fill_sram_inverted $T=3162 1306 1 0 $X=3138 $Y=590
XX73A2B17220_19 GND! VDD! 127 159 fill_sram_inverted $T=3330 1306 1 0 $X=3306 $Y=590
XX73A2B17239_1 GND! VDD! 126 160 fill_sram_inverted $T=306 13078 1 0 $X=282 $Y=12362
XX73A2B17239_2 GND! VDD! 126 160 fill_sram_inverted $T=474 13078 1 0 $X=450 $Y=12362
XX73A2B17239_3 GND! VDD! 126 160 fill_sram_inverted $T=642 13078 1 0 $X=618 $Y=12362
XX73A2B17239_4 GND! VDD! 126 160 fill_sram_inverted $T=810 13078 1 0 $X=786 $Y=12362
XX73A2B17239_5 GND! VDD! 126 160 fill_sram_inverted $T=978 13078 1 0 $X=954 $Y=12362
XX73A2B17239_6 GND! VDD! 126 160 fill_sram_inverted $T=1146 13078 1 0 $X=1122 $Y=12362
XX73A2B17239_7 GND! VDD! 126 160 fill_sram_inverted $T=1314 13078 1 0 $X=1290 $Y=12362
XX73A2B17239_8 GND! VDD! 126 160 fill_sram_inverted $T=1482 13078 1 0 $X=1458 $Y=12362
XX73A2B17239_9 GND! VDD! 126 160 fill_sram_inverted $T=1650 13078 1 0 $X=1626 $Y=12362
XX73A2B17239_10 GND! VDD! 126 160 fill_sram_inverted $T=1818 13078 1 0 $X=1794 $Y=12362
XX73A2B17239_11 GND! VDD! 126 160 fill_sram_inverted $T=1986 13078 1 0 $X=1962 $Y=12362
XX73A2B17239_12 GND! VDD! 126 160 fill_sram_inverted $T=2154 13078 1 0 $X=2130 $Y=12362
XX73A2B17239_13 GND! VDD! 126 160 fill_sram_inverted $T=2322 13078 1 0 $X=2298 $Y=12362
XX73A2B17239_14 GND! VDD! 126 160 fill_sram_inverted $T=2490 13078 1 0 $X=2466 $Y=12362
XX73A2B17239_15 GND! VDD! 126 160 fill_sram_inverted $T=2658 13078 1 0 $X=2634 $Y=12362
XX73A2B17239_16 GND! VDD! 126 160 fill_sram_inverted $T=2826 13078 1 0 $X=2802 $Y=12362
XX73A2B17239_17 GND! VDD! 126 160 fill_sram_inverted $T=2994 13078 1 0 $X=2970 $Y=12362
XX73A2B17239_18 GND! VDD! 126 160 fill_sram_inverted $T=3162 13078 1 0 $X=3138 $Y=12362
XX73A2B17239_19 GND! VDD! 126 160 fill_sram_inverted $T=3330 13078 1 0 $X=3306 $Y=12362
XX73A2B17239_20 GND! VDD! 126 160 fill_sram_inverted $T=3498 13078 1 0 $X=3474 $Y=12362
XX73A2B17239_21 GND! VDD! 126 160 fill_sram_inverted $T=3666 13078 1 0 $X=3642 $Y=12362
XX73A2B17239_22 GND! VDD! 126 160 fill_sram_inverted $T=3834 13078 1 0 $X=3810 $Y=12362
XX73A2B17261_1 GND! VDD! 128 158 fill_sram_inverted $T=306 14386 1 0 $X=282 $Y=13670
XX73A2B17261_2 GND! VDD! 128 158 fill_sram_inverted $T=474 14386 1 0 $X=450 $Y=13670
XX73A2B17261_3 GND! VDD! 128 158 fill_sram_inverted $T=642 14386 1 0 $X=618 $Y=13670
XX73A2B17261_4 GND! VDD! 128 158 fill_sram_inverted $T=810 14386 1 0 $X=786 $Y=13670
XX73A2B17261_5 GND! VDD! 128 158 fill_sram_inverted $T=978 14386 1 0 $X=954 $Y=13670
XX73A2B17261_6 GND! VDD! 128 158 fill_sram_inverted $T=1146 14386 1 0 $X=1122 $Y=13670
XX73A2B17261_7 GND! VDD! 128 158 fill_sram_inverted $T=1314 14386 1 0 $X=1290 $Y=13670
XX73A2B17261_8 GND! VDD! 128 158 fill_sram_inverted $T=1482 14386 1 0 $X=1458 $Y=13670
XX73A2B17261_9 GND! VDD! 128 158 fill_sram_inverted $T=1650 14386 1 0 $X=1626 $Y=13670
XX73A2B17261_10 GND! VDD! 128 158 fill_sram_inverted $T=1818 14386 1 0 $X=1794 $Y=13670
XX73A2B17261_11 GND! VDD! 128 158 fill_sram_inverted $T=1986 14386 1 0 $X=1962 $Y=13670
XX73A2B17261_12 GND! VDD! 128 158 fill_sram_inverted $T=2154 14386 1 0 $X=2130 $Y=13670
XX73A2B17261_13 GND! VDD! 128 158 fill_sram_inverted $T=2322 14386 1 0 $X=2298 $Y=13670
XX73A2B17261_14 GND! VDD! 128 158 fill_sram_inverted $T=2490 14386 1 0 $X=2466 $Y=13670
XX73A2B17261_15 GND! VDD! 128 158 fill_sram_inverted $T=2658 14386 1 0 $X=2634 $Y=13670
XX73A2B17261_16 GND! VDD! 128 158 fill_sram_inverted $T=2826 14386 1 0 $X=2802 $Y=13670
XX73A2B17261_17 GND! VDD! 128 158 fill_sram_inverted $T=2994 14386 1 0 $X=2970 $Y=13670
XX73A2B17261_18 GND! VDD! 128 158 fill_sram_inverted $T=3162 14386 1 0 $X=3138 $Y=13670
XX73A2B17261_19 GND! VDD! 128 158 fill_sram_inverted $T=3330 14386 1 0 $X=3306 $Y=13670
XX73A2B17280 57 69 43 GND! VDD! 129 161 buffer_top $T=2970 6470 0 0 $X=2970 $Y=6476
XX73A2B17281 55 70 42 GND! VDD! 130 162 buffer_top $T=2970 5162 0 0 $X=2970 $Y=5168
XX73A2B17282 53 71 38 GND! VDD! 131 163 buffer_top $T=2970 3854 0 0 $X=2970 $Y=3860
XX73A2B17283 51 72 37 GND! VDD! 132 164 buffer_top $T=2970 2546 0 0 $X=2970 $Y=2552
XX73A2B17284 49 73 36 GND! VDD! 127 165 buffer_top $T=2970 1238 0 0 $X=2970 $Y=1244
XX73A2B17285 59 74 44 GND! VDD! 133 166 buffer_top $T=2970 7778 0 0 $X=2970 $Y=7784
XX73A2B17286 61 75 47 GND! VDD! 134 167 buffer_top $T=2970 9086 0 0 $X=2970 $Y=9092
XX73A2B17287 63 76 48 GND! VDD! 135 168 buffer_top $T=2970 10394 0 0 $X=2970 $Y=10400
XX73A2B17288 A<4> 77 142 143 144 145 147 146 149 148 WENB 
+	16 22 18 23 17 10 21 12 9 15 19 
+	11 20 24 13 14 D<0> D<1> D<2> D<3> GND! VDD! 
+	VDD! GND! 128 126 136 169 158 column_decoder_write $T=3528 13010 0 0 $X=3474 $Y=13016
XX73A2B17289_1 GND! VDD! 137 160 fill_sram $T=2994 11772 0 0 $X=2970 $Y=11708
XX73A2B17289_2 GND! VDD! 137 160 fill_sram $T=3162 11772 0 0 $X=3138 $Y=11708
XX73A2B17289_3 GND! VDD! 137 160 fill_sram $T=3330 11772 0 0 $X=3306 $Y=11708
XX73A2B17289_4 GND! VDD! 137 160 fill_sram $T=3498 11772 0 0 $X=3474 $Y=11708
XX73A2B17289_5 GND! VDD! 137 160 fill_sram $T=3666 11772 0 0 $X=3642 $Y=11708
XX73A2B17289_6 GND! VDD! 137 160 fill_sram $T=3834 11772 0 0 $X=3810 $Y=11708
XX73A2B17295_1 GND! VDD! 128 169 fill_sram $T=306 14388 0 0 $X=282 $Y=14324
XX73A2B17295_2 GND! VDD! 128 169 fill_sram $T=474 14388 0 0 $X=450 $Y=14324
XX73A2B17295_3 GND! VDD! 128 169 fill_sram $T=642 14388 0 0 $X=618 $Y=14324
XX73A2B17295_4 GND! VDD! 128 169 fill_sram $T=810 14388 0 0 $X=786 $Y=14324
XX73A2B17295_5 GND! VDD! 128 169 fill_sram $T=978 14388 0 0 $X=954 $Y=14324
XX73A2B17295_6 GND! VDD! 128 169 fill_sram $T=1146 14388 0 0 $X=1122 $Y=14324
XX73A2B17295_7 GND! VDD! 128 169 fill_sram $T=1314 14388 0 0 $X=1290 $Y=14324
XX73A2B17295_8 GND! VDD! 128 169 fill_sram $T=1482 14388 0 0 $X=1458 $Y=14324
XX73A2B17295_9 GND! VDD! 128 169 fill_sram $T=1650 14388 0 0 $X=1626 $Y=14324
XX73A2B17295_10 GND! VDD! 128 169 fill_sram $T=1818 14388 0 0 $X=1794 $Y=14324
XX73A2B17295_11 GND! VDD! 128 169 fill_sram $T=1986 14388 0 0 $X=1962 $Y=14324
XX73A2B17295_12 GND! VDD! 128 169 fill_sram $T=2154 14388 0 0 $X=2130 $Y=14324
XX73A2B17295_13 GND! VDD! 128 169 fill_sram $T=2322 14388 0 0 $X=2298 $Y=14324
XX73A2B17295_14 GND! VDD! 128 169 fill_sram $T=2490 14388 0 0 $X=2466 $Y=14324
XX73A2B17295_15 GND! VDD! 128 169 fill_sram $T=2658 14388 0 0 $X=2634 $Y=14324
XX73A2B17295_16 GND! VDD! 128 169 fill_sram $T=2826 14388 0 0 $X=2802 $Y=14324
XX73A2B17295_17 GND! VDD! 128 169 fill_sram $T=2994 14388 0 0 $X=2970 $Y=14324
XX73A2B17295_18 GND! VDD! 128 169 fill_sram $T=3162 14388 0 0 $X=3138 $Y=14324
XX73A2B17295_19 GND! VDD! 128 169 fill_sram $T=3330 14388 0 0 $X=3306 $Y=14324
XX73A2B172114_1 GND! VDD! 138 159 fill_sram $T=306 0 0 0 $X=282 $Y=-64
XX73A2B172114_2 GND! VDD! 138 159 fill_sram $T=474 0 0 0 $X=450 $Y=-64
XX73A2B172114_3 GND! VDD! 138 159 fill_sram $T=642 0 0 0 $X=618 $Y=-64
XX73A2B172114_4 GND! VDD! 138 159 fill_sram $T=810 0 0 0 $X=786 $Y=-64
XX73A2B172114_5 GND! VDD! 138 159 fill_sram $T=978 0 0 0 $X=954 $Y=-64
XX73A2B172114_6 GND! VDD! 138 159 fill_sram $T=1146 0 0 0 $X=1122 $Y=-64
XX73A2B172114_7 GND! VDD! 138 159 fill_sram $T=1314 0 0 0 $X=1290 $Y=-64
XX73A2B172114_8 GND! VDD! 138 159 fill_sram $T=1482 0 0 0 $X=1458 $Y=-64
XX73A2B172114_9 GND! VDD! 138 159 fill_sram $T=1650 0 0 0 $X=1626 $Y=-64
XX73A2B172114_10 GND! VDD! 138 159 fill_sram $T=1818 0 0 0 $X=1794 $Y=-64
XX73A2B172114_11 GND! VDD! 138 159 fill_sram $T=1986 0 0 0 $X=1962 $Y=-64
XX73A2B172114_12 GND! VDD! 138 159 fill_sram $T=2154 0 0 0 $X=2130 $Y=-64
XX73A2B172114_13 GND! VDD! 138 159 fill_sram $T=2322 0 0 0 $X=2298 $Y=-64
XX73A2B172114_14 GND! VDD! 138 159 fill_sram $T=2490 0 0 0 $X=2466 $Y=-64
XX73A2B172114_15 GND! VDD! 138 159 fill_sram $T=2658 0 0 0 $X=2634 $Y=-64
XX73A2B172114_16 GND! VDD! 138 159 fill_sram $T=2826 0 0 0 $X=2802 $Y=-64
XX73A2B172114_17 GND! VDD! 138 159 fill_sram $T=2994 0 0 0 $X=2970 $Y=-64
XX73A2B172114_18 GND! VDD! 138 159 fill_sram $T=3162 0 0 0 $X=3138 $Y=-64
XX73A2B172114_19 GND! VDD! 138 159 fill_sram $T=3330 0 0 0 $X=3306 $Y=-64
XX73A2B172114_20 GND! VDD! 138 159 fill_sram $T=3498 0 0 0 $X=3474 $Y=-64
XX73A2B172114_21 GND! VDD! 138 159 fill_sram $T=3666 0 0 0 $X=3642 $Y=-64
XX73A2B172114_22 GND! VDD! 138 159 fill_sram $T=3834 0 0 0 $X=3810 $Y=-64
XX73A2B172114_23 GND! VDD! 138 159 fill_sram $T=4002 0 0 0 $X=3977 $Y=-64
XX73A2B172114_24 GND! VDD! 138 159 fill_sram $T=4170 0 0 0 $X=4146 $Y=-64
XX73A2B172114_25 GND! VDD! 138 159 fill_sram $T=4338 0 0 0 $X=4314 $Y=-64
XX73A2B172114_26 GND! VDD! 138 159 fill_sram $T=4506 0 0 0 $X=4482 $Y=-64
XX73A2B172140 58 78 40 GND! VDD! 133 161 buffer_top_inverted $T=2970 7916 1 0 $X=2970 $Y=7130
XX73A2B172141 56 79 39 GND! VDD! 129 162 buffer_top_inverted $T=2970 6608 1 0 $X=2970 $Y=5822
XX73A2B172142 54 80 35 GND! VDD! 130 163 buffer_top_inverted $T=2970 5300 1 0 $X=2970 $Y=4513
XX73A2B172143 52 81 34 GND! VDD! 131 164 buffer_top_inverted $T=2970 3992 1 0 $X=2970 $Y=3206
XX73A2B172144 50 82 33 GND! VDD! 132 165 buffer_top_inverted $T=2970 2684 1 0 $X=2970 $Y=1898
XX73A2B172145 60 83 41 GND! VDD! 134 166 buffer_top_inverted $T=2970 9224 1 0 $X=2970 $Y=8438
XX73A2B172146 62 84 45 GND! VDD! 135 167 buffer_top_inverted $T=2970 10532 1 0 $X=2970 $Y=9746
XX73A2B172147 64 85 46 GND! VDD! 137 168 buffer_top_inverted $T=2970 11840 1 0 $X=2970 $Y=11054
XX73A2B172148 CLK 16 17 18 19 20 13 21 9 22 10 
+	23 11 24 14 12 15 GND! VDD! GND! 137 126 
+	160 bitline_conditioning $T=4032 11772 0 0 $X=3978 $Y=11708
XX73A2B172149 CLK A<1> A<0> A<2> A<3> 86 139 141 140 33 34 
+	35 36 37 38 39 40 41 42 43 44 45 
+	46 47 48 GND! GND! VDD! GND! VDD! GND! VDD! GND! 
+	VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 132 
+	131 127 130 129 133 134 135 137 165 164 163 
+	162 161 166 167 168 160 row_decoder_4_16 $T=336 1308 0 0 $X=282 $Y=1244
XX73A2B172150 A<4> 87 9 15 WENB 68 13 14 67 19 11 
+	66 17 10 65 VDD! GND! 127 159 150 151 152 
+	153 154 155 156 157 column_decoder_read $T=2966 590 0 0 $X=3474 $Y=590
XX73A2B172151 16 17 18 19 20 13 21 9 22 10 23 
+	11 24 14 12 15 52 50 51 49 56 54 
+	55 53 60 58 59 57 64 62 63 61 VDD! 
+	GND! VDD! GND! VDD! GND! GND! VDD! VDD! GND! GND! VDD! 
+	GND! VDD! GND! VDD! GND! 88 89 90 91 92 93 
+	94 95 96 97 98 99 100 101 102 103 104 
+	105 106 107 108 109 110 111 112 113 114 115 
+	116 117 118 119 133 134 137 135 130 129 131 
+	132 127 161 166 168 167 163 162 164 165 sram_array_16r_8c $T=4032 1308 0 0 $X=3978 $Y=1244
XX73A2B172152 VDD! GND! 126 137 128 133 135 134 127 132 131 
+	130 129 138 136 158 168 160 161 167 166 159 
+	165 164 163 162 169 sram_lvs_grid $T=-46 -70 0 0 $X=-54 $Y=-64
XX73A2B172153 VDD! GND! 126 137 128 133 135 134 127 132 131 
+	130 129 138 136 158 168 160 161 167 166 159 
+	165 164 163 162 169 sram_lvs_grid $T=11882 -70 0 0 $X=11874 $Y=-64
XX73A2B172154 120 68 121 67 122 66 123 65 GND! VDD! Q<0> 
+	Q<1> Q<2> Q<3> 138 159 buffer_array $T=4650 -70 0 0 $X=4650 $Y=-64
.ends top_level
