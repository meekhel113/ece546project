*  Generated for: PrimeSim
*  Design library name: project_backup
*  Design cell name: top_level_tb
*  Design view name: schematic
.option search='/afs/eos.ncsu.edu/lockers/research/ece/wdavis/tech/FreePDK3/hspice/models'

.param clkperiod=0.21n clkrise=5p vdd=0.8
.option PARHIER = LOCAL
.option PORT_VOLTAGE_SCALE_TO_2X = 1

.option WDF=1
.temp 25
.lib 'fet.mod' nfet_typ
.lib 'fet.mod' pfet_typ
.vec '/afs/unity.ncsu.edu/users/s/ssjoseph/ECE546/PROJECT/ece546project/invec_local.dat'

.vec '/afs/unity.ncsu.edu/users/s/ssjoseph/ECE546/PROJECT/ece546project/outvec_local.dat'


*Custom Compiler Version S-2021.09
*Thu Apr 21 18:04:47 2022

.global 0 gnd! vdd!
********************************************************************************
* Library          : project_backup
* Cell             : inputbuf
* View             : schematic
* View Search List : starrc hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt inputbuf out in
m11 out net7 vdd! pfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
m10 net7 in vdd! pfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
m9 out net7 gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m8 net7 in gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
.ends inputbuf

********************************************************************************
* Library          : project_backup
* Cell             : top_level
* View             : starrc
* View Search List : starrc hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt top_level a<0> a<1> a<2> a<3> a<4> clk d<0> d<1> d<2> d<3> q<0> q<1>
+ q<2> q<3> wenb
mi11|m124 net266 a<0> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m181 net266 i11|net698 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m167 net266 i11|net699 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m153 net266 i11|net700 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m126 net282 a<0> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m183 net282 i11|net698 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m100 net282 a<2> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m157 net282 i11|net700 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m128 net286 a<0> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m185 net286 i11|net698 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m171 net286 i11|net699 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m88 net286 a<3> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m130 net290 a<0> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m187 net290 i11|net698 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m105 net290 a<2> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m92 net290 a<3> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m195 net265 i11|net697 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m180 net265 i11|net698 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m166 net265 i11|net699 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m152 net265 i11|net700 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m193 net281 i11|net697 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m182 net281 i11|net698 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m99 net281 a<2> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m156 net281 i11|net700 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m191 net285 i11|net697 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m184 net285 i11|net698 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m170 net285 i11|net699 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m87 net285 a<3> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m189 net289 i11|net697 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m186 net289 i11|net698 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m106 net289 a<2> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m91 net289 a<3> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|i234|m0@2 gnd! a<2> i11|net699 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi11|m173 net288 i11|net699 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m102 net284 a<2> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m169 net268 i11|net699 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|i235|m0 i11|net700 a<3> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi11|m90 net288 a<3> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m190 net287 i11|net697 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m192 net283 i11|net697 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m194 net267 i11|net697 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m159 net284 i11|net700 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|i232|m0 i11|net697 a<0> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi11|i232|m0@2 gnd! a<0> i11|net697 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi11|m119 net287 a<1> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m115 net283 a<1> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m111 net267 a<1> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m172 net287 i11|net699 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m101 net283 a<2> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m168 net267 i11|net699 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|i233|m0 i11|net698 a<1> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi11|i233|m0@2 gnd! a<1> i11|net698 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi11|m155 net268 i11|net700 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m89 net287 a<3> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m158 net283 i11|net700 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m154 net267 i11|net700 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi11|m129 net288 a<0> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m127 net284 a<0> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m125 net268 a<0> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|i234|m0 i11|net699 a<2> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi11|m118 net288 a<1> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m114 net284 a<1> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m112 net268 a<1> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|i235|m0@2 gnd! a<3> i11|net700 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi40|i1|i1|m0@2 gnd! i40|i1|net4 q<2> nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi40|i2|i0|m0 i40|i2|net4 net225 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi40|i2|i0|m0@2 gnd! net225 i40|i2|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi40|i2|i1|m0 q<1> i40|i2|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi40|i2|i1|m0@2 gnd! i40|i2|net4 q<1> nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi40|i3|i0|m0 i40|i3|net4 net355 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi40|i3|i0|m0@2 gnd! net355 i40|i3|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi40|i3|i1|m0 q<0> i40|i3|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi40|i0|i0|m0 i40|i0|net4 net229 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi40|i0|i0|m0@2 gnd! net229 i40|i0|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi40|i0|i1|m0 q<3> i40|i0|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi40|i0|i1|m0@2 gnd! i40|i0|net4 q<3> nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi40|i1|i0|m0 i40|i1|net4 net227 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi40|i1|i0|m0@2 gnd! net227 i40|i1|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi40|i1|i1|m0 q<2> i40|i1|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi40|i3|i1|m0@2 gnd! i40|i3|net4 q<0> nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i59|i1|m11 bl<1> net262 i0|i59|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i57|i0|m10 blb<0> net263 i0|i57|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i59|i0|m10 blb<0> net262 i0|i59|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i57|i0|m1 gnd! i0|i57|i0|q i0|i57|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i59|i0|m1 gnd! i0|i59|i0|q i0|i59|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i57|i0|m3 i0|i57|i0|q i0|i57|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i57|i3|m10 blb<3> net263 i0|i57|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i59|i3|m10 blb<3> net262 i0|i59|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i57|i3|m1 gnd! i0|i57|i3|q i0|i57|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i59|i0|m3 i0|i59|i0|q i0|i59|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i59|i3|m1 gnd! i0|i59|i3|q i0|i59|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i57|i3|m3 i0|i57|i3|q i0|i57|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i59|i3|m3 i0|i59|i3|q i0|i59|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i57|i3|m11 bl<3> net263 i0|i57|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i59|i3|m11 bl<3> net262 i0|i59|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i57|i2|m10 blb<2> net263 i0|i57|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i59|i2|m10 blb<2> net262 i0|i59|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i57|i2|m1 gnd! i0|i57|i2|q i0|i57|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i59|i2|m1 gnd! i0|i59|i2|q i0|i59|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i57|i2|m3 i0|i57|i2|q i0|i57|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i57|i0|m11 bl<0> net263 i0|i57|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i59|i2|m3 i0|i59|i2|q i0|i59|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i57|i2|m11 bl<2> net263 i0|i57|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i59|i2|m11 bl<2> net262 i0|i59|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i57|i1|m10 blb<1> net263 i0|i57|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i59|i1|m10 blb<1> net262 i0|i59|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i57|i1|m1 gnd! i0|i57|i1|q i0|i57|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i59|i1|m1 gnd! i0|i59|i1|q i0|i59|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i57|i1|m3 i0|i57|i1|q i0|i57|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i59|i1|m3 i0|i59|i1|q i0|i59|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i57|i1|m11 bl<1> net263 i0|i57|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i59|i0|m11 bl<0> net262 i0|i59|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i51|i1|m11 bl<1> net270 i0|i51|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i49|i0|m10 blb<0> net271 i0|i49|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i51|i0|m10 blb<0> net270 i0|i51|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i49|i0|m1 gnd! i0|i49|i0|q i0|i49|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i51|i0|m1 gnd! i0|i51|i0|q i0|i51|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i49|i0|m3 i0|i49|i0|q i0|i49|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i49|i3|m10 blb<3> net271 i0|i49|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i51|i3|m10 blb<3> net270 i0|i51|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i49|i3|m1 gnd! i0|i49|i3|q i0|i49|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i51|i0|m3 i0|i51|i0|q i0|i51|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i51|i3|m1 gnd! i0|i51|i3|q i0|i51|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i49|i3|m3 i0|i49|i3|q i0|i49|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i51|i3|m3 i0|i51|i3|q i0|i51|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i49|i3|m11 bl<3> net271 i0|i49|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i51|i3|m11 bl<3> net270 i0|i51|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i49|i2|m10 blb<2> net271 i0|i49|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i51|i2|m10 blb<2> net270 i0|i51|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i49|i2|m1 gnd! i0|i49|i2|q i0|i49|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i51|i2|m1 gnd! i0|i51|i2|q i0|i51|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i49|i2|m3 i0|i49|i2|q i0|i49|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i49|i0|m11 bl<0> net271 i0|i49|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i51|i2|m3 i0|i51|i2|q i0|i51|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i49|i2|m11 bl<2> net271 i0|i49|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i51|i2|m11 bl<2> net270 i0|i51|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i49|i1|m10 blb<1> net271 i0|i49|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i51|i1|m10 blb<1> net270 i0|i51|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i49|i1|m1 gnd! i0|i49|i1|q i0|i49|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i51|i1|m1 gnd! i0|i51|i1|q i0|i51|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i49|i1|m3 i0|i49|i1|q i0|i49|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i51|i1|m3 i0|i51|i1|q i0|i51|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i49|i1|m11 bl<1> net271 i0|i49|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i51|i0|m11 bl<0> net270 i0|i51|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i43|i1|m11 bl<1> net274 i0|i43|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i41|i0|m10 blb<0> net275 i0|i41|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i43|i0|m10 blb<0> net274 i0|i43|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i41|i0|m1 gnd! i0|i41|i0|q i0|i41|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i43|i0|m1 gnd! i0|i43|i0|q i0|i43|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i41|i0|m3 i0|i41|i0|q i0|i41|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i41|i3|m10 blb<3> net275 i0|i41|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i43|i3|m10 blb<3> net274 i0|i43|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i41|i3|m1 gnd! i0|i41|i3|q i0|i41|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i43|i0|m3 i0|i43|i0|q i0|i43|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i43|i3|m1 gnd! i0|i43|i3|q i0|i43|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i41|i3|m3 i0|i41|i3|q i0|i41|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i43|i3|m3 i0|i43|i3|q i0|i43|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i41|i3|m11 bl<3> net275 i0|i41|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i43|i3|m11 bl<3> net274 i0|i43|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i41|i2|m10 blb<2> net275 i0|i41|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i43|i2|m10 blb<2> net274 i0|i43|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i41|i2|m1 gnd! i0|i41|i2|q i0|i41|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i43|i2|m1 gnd! i0|i43|i2|q i0|i43|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i41|i2|m3 i0|i41|i2|q i0|i41|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i41|i0|m11 bl<0> net275 i0|i41|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i43|i2|m3 i0|i43|i2|q i0|i43|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i41|i2|m11 bl<2> net275 i0|i41|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i43|i2|m11 bl<2> net274 i0|i43|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i41|i1|m10 blb<1> net275 i0|i41|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i43|i1|m10 blb<1> net274 i0|i43|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i41|i1|m1 gnd! i0|i41|i1|q i0|i41|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i43|i1|m1 gnd! i0|i43|i1|q i0|i43|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i41|i1|m3 i0|i41|i1|q i0|i41|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i43|i1|m3 i0|i43|i1|q i0|i43|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i41|i1|m11 bl<1> net275 i0|i41|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i43|i0|m11 bl<0> net274 i0|i43|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i35|i1|m11 bl<1> net278 i0|i35|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i33|i0|m10 blb<0> net279 i0|i33|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i35|i0|m10 blb<0> net278 i0|i35|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i33|i0|m1 gnd! i0|i33|i0|q i0|i33|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i35|i0|m1 gnd! i0|i35|i0|q i0|i35|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i33|i0|m3 i0|i33|i0|q i0|i33|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i33|i3|m10 blb<3> net279 i0|i33|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i35|i3|m10 blb<3> net278 i0|i35|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i33|i3|m1 gnd! i0|i33|i3|q i0|i33|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i35|i0|m3 i0|i35|i0|q i0|i35|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i35|i3|m1 gnd! i0|i35|i3|q i0|i35|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i33|i3|m3 i0|i33|i3|q i0|i33|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i35|i3|m3 i0|i35|i3|q i0|i35|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i33|i3|m11 bl<3> net279 i0|i33|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i35|i3|m11 bl<3> net278 i0|i35|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i33|i2|m10 blb<2> net279 i0|i33|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i35|i2|m10 blb<2> net278 i0|i35|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i33|i2|m1 gnd! i0|i33|i2|q i0|i33|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i35|i2|m1 gnd! i0|i35|i2|q i0|i35|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i33|i2|m3 i0|i33|i2|q i0|i33|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i33|i0|m11 bl<0> net279 i0|i33|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i35|i2|m3 i0|i35|i2|q i0|i35|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i33|i2|m11 bl<2> net279 i0|i33|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i35|i2|m11 bl<2> net278 i0|i35|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i33|i1|m10 blb<1> net279 i0|i33|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i35|i1|m10 blb<1> net278 i0|i35|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i33|i1|m1 gnd! i0|i33|i1|q i0|i33|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i35|i1|m1 gnd! i0|i35|i1|q i0|i35|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i33|i1|m3 i0|i33|i1|q i0|i33|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i35|i1|m3 i0|i35|i1|q i0|i35|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i33|i1|m11 bl<1> net279 i0|i33|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i35|i0|m11 bl<0> net278 i0|i35|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i58|i1|m11 bl<5> net262 i0|i58|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i56|i0|m10 blb<4> net263 i0|i56|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i58|i0|m10 blb<4> net262 i0|i58|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i56|i0|m1 gnd! i0|i56|i0|q i0|i56|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i58|i0|m1 gnd! i0|i58|i0|q i0|i58|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i56|i0|m3 i0|i56|i0|q i0|i56|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i56|i3|m10 blb<7> net263 i0|i56|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i58|i3|m10 blb<7> net262 i0|i58|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i56|i3|m1 gnd! i0|i56|i3|q i0|i56|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i58|i0|m3 i0|i58|i0|q i0|i58|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i58|i3|m1 gnd! i0|i58|i3|q i0|i58|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i56|i3|m3 i0|i56|i3|q i0|i56|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i58|i3|m3 i0|i58|i3|q i0|i58|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i56|i3|m11 bl<7> net263 i0|i56|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i58|i3|m11 bl<7> net262 i0|i58|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i56|i2|m10 blb<6> net263 i0|i56|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i58|i2|m10 blb<6> net262 i0|i58|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i56|i2|m1 gnd! i0|i56|i2|q i0|i56|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i58|i2|m1 gnd! i0|i58|i2|q i0|i58|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i56|i2|m3 i0|i56|i2|q i0|i56|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i56|i0|m11 bl<4> net263 i0|i56|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i58|i2|m3 i0|i58|i2|q i0|i58|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i56|i2|m11 bl<6> net263 i0|i56|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i58|i2|m11 bl<6> net262 i0|i58|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i56|i1|m10 blb<5> net263 i0|i56|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i58|i1|m10 blb<5> net262 i0|i58|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i56|i1|m1 gnd! i0|i56|i1|q i0|i56|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i58|i1|m1 gnd! i0|i58|i1|q i0|i58|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i56|i1|m3 i0|i56|i1|q i0|i56|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i58|i1|m3 i0|i58|i1|q i0|i58|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i56|i1|m11 bl<5> net263 i0|i56|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i58|i0|m11 bl<4> net262 i0|i58|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i50|i1|m11 bl<5> net270 i0|i50|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i48|i0|m10 blb<4> net271 i0|i48|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i50|i0|m10 blb<4> net270 i0|i50|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i48|i0|m1 gnd! i0|i48|i0|q i0|i48|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i50|i0|m1 gnd! i0|i50|i0|q i0|i50|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i48|i0|m3 i0|i48|i0|q i0|i48|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i48|i3|m10 blb<7> net271 i0|i48|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i50|i3|m10 blb<7> net270 i0|i50|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i48|i3|m1 gnd! i0|i48|i3|q i0|i48|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i50|i0|m3 i0|i50|i0|q i0|i50|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i50|i3|m1 gnd! i0|i50|i3|q i0|i50|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i48|i3|m3 i0|i48|i3|q i0|i48|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i50|i3|m3 i0|i50|i3|q i0|i50|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i48|i3|m11 bl<7> net271 i0|i48|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i50|i3|m11 bl<7> net270 i0|i50|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i48|i2|m10 blb<6> net271 i0|i48|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i50|i2|m10 blb<6> net270 i0|i50|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i48|i2|m1 gnd! i0|i48|i2|q i0|i48|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i50|i2|m1 gnd! i0|i50|i2|q i0|i50|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i48|i2|m3 i0|i48|i2|q i0|i48|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i48|i0|m11 bl<4> net271 i0|i48|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i50|i2|m3 i0|i50|i2|q i0|i50|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i48|i2|m11 bl<6> net271 i0|i48|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i50|i2|m11 bl<6> net270 i0|i50|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i48|i1|m10 blb<5> net271 i0|i48|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i50|i1|m10 blb<5> net270 i0|i50|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i48|i1|m1 gnd! i0|i48|i1|q i0|i48|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i50|i1|m1 gnd! i0|i50|i1|q i0|i50|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i48|i1|m3 i0|i48|i1|q i0|i48|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i50|i1|m3 i0|i50|i1|q i0|i50|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i48|i1|m11 bl<5> net271 i0|i48|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i50|i0|m11 bl<4> net270 i0|i50|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i42|i1|m11 bl<5> net274 i0|i42|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i40|i0|m10 blb<4> net275 i0|i40|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i42|i0|m10 blb<4> net274 i0|i42|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i40|i0|m1 gnd! i0|i40|i0|q i0|i40|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i42|i0|m1 gnd! i0|i42|i0|q i0|i42|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i40|i0|m3 i0|i40|i0|q i0|i40|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i40|i3|m10 blb<7> net275 i0|i40|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i42|i3|m10 blb<7> net274 i0|i42|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i40|i3|m1 gnd! i0|i40|i3|q i0|i40|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i42|i0|m3 i0|i42|i0|q i0|i42|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i42|i3|m1 gnd! i0|i42|i3|q i0|i42|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i40|i3|m3 i0|i40|i3|q i0|i40|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i42|i3|m3 i0|i42|i3|q i0|i42|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i40|i3|m11 bl<7> net275 i0|i40|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i42|i3|m11 bl<7> net274 i0|i42|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i40|i2|m10 blb<6> net275 i0|i40|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i42|i2|m10 blb<6> net274 i0|i42|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i40|i2|m1 gnd! i0|i40|i2|q i0|i40|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i42|i2|m1 gnd! i0|i42|i2|q i0|i42|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i40|i2|m3 i0|i40|i2|q i0|i40|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i40|i0|m11 bl<4> net275 i0|i40|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i42|i2|m3 i0|i42|i2|q i0|i42|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i40|i2|m11 bl<6> net275 i0|i40|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i42|i2|m11 bl<6> net274 i0|i42|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i40|i1|m10 blb<5> net275 i0|i40|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i42|i1|m10 blb<5> net274 i0|i42|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i40|i1|m1 gnd! i0|i40|i1|q i0|i40|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i42|i1|m1 gnd! i0|i42|i1|q i0|i42|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i40|i1|m3 i0|i40|i1|q i0|i40|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i42|i1|m3 i0|i42|i1|q i0|i42|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i40|i1|m11 bl<5> net275 i0|i40|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i42|i0|m11 bl<4> net274 i0|i42|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i34|i1|m11 bl<5> net278 i0|i34|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i32|i0|m10 blb<4> net279 i0|i32|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i34|i0|m10 blb<4> net278 i0|i34|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i32|i0|m1 gnd! i0|i32|i0|q i0|i32|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i34|i0|m1 gnd! i0|i34|i0|q i0|i34|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i32|i0|m3 i0|i32|i0|q i0|i32|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i32|i3|m10 blb<7> net279 i0|i32|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i34|i3|m10 blb<7> net278 i0|i34|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i32|i3|m1 gnd! i0|i32|i3|q i0|i32|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i34|i0|m3 i0|i34|i0|q i0|i34|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i34|i3|m1 gnd! i0|i34|i3|q i0|i34|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i32|i3|m3 i0|i32|i3|q i0|i32|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i34|i3|m3 i0|i34|i3|q i0|i34|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i32|i3|m11 bl<7> net279 i0|i32|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i34|i3|m11 bl<7> net278 i0|i34|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i32|i2|m10 blb<6> net279 i0|i32|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i34|i2|m10 blb<6> net278 i0|i34|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i32|i2|m1 gnd! i0|i32|i2|q i0|i32|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i34|i2|m1 gnd! i0|i34|i2|q i0|i34|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i32|i2|m3 i0|i32|i2|q i0|i32|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i32|i0|m11 bl<4> net279 i0|i32|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i34|i2|m3 i0|i34|i2|q i0|i34|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i32|i2|m11 bl<6> net279 i0|i32|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i34|i2|m11 bl<6> net278 i0|i34|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i32|i1|m10 blb<5> net279 i0|i32|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i34|i1|m10 blb<5> net278 i0|i34|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i32|i1|m1 gnd! i0|i32|i1|q i0|i32|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i34|i1|m1 gnd! i0|i34|i1|q i0|i34|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i32|i1|m3 i0|i32|i1|q i0|i32|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i34|i1|m3 i0|i34|i1|q i0|i34|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i32|i1|m11 bl<5> net279 i0|i32|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i34|i0|m11 bl<4> net278 i0|i34|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i46|i2|m11 bl<6> net272 i0|i46|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i52|i2|m11 bl<6> net269 i0|i52|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i54|i2|m11 bl<6> net264 i0|i54|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i44|i1|m10 blb<5> net273 i0|i44|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i46|i1|m10 blb<5> net272 i0|i46|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i52|i1|m10 blb<5> net269 i0|i52|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i54|i1|m10 blb<5> net264 i0|i54|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i44|i1|m1 gnd! i0|i44|i1|q i0|i44|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i46|i1|m1 gnd! i0|i46|i1|q i0|i46|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i52|i1|m1 gnd! i0|i52|i1|q i0|i52|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i55|i0|m1 gnd! i0|i55|i0|q i0|i55|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i54|i1|m1 gnd! i0|i54|i1|q i0|i54|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i44|i1|m3 i0|i44|i1|q i0|i44|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i46|i1|m3 i0|i46|i1|q i0|i46|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i52|i1|m3 i0|i52|i1|q i0|i52|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i54|i1|m3 i0|i54|i1|q i0|i54|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i44|i1|m11 bl<5> net273 i0|i44|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i46|i1|m11 bl<5> net272 i0|i46|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i52|i1|m11 bl<5> net269 i0|i52|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i54|i1|m11 bl<5> net264 i0|i54|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i44|i0|m10 blb<4> net273 i0|i44|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i45|i0|m3 i0|i45|i0|q i0|i45|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i46|i0|m10 blb<4> net272 i0|i46|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i52|i0|m10 blb<4> net269 i0|i52|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i54|i0|m10 blb<4> net264 i0|i54|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i44|i0|m1 gnd! i0|i44|i0|q i0|i44|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i46|i0|m1 gnd! i0|i46|i0|q i0|i46|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i52|i0|m1 gnd! i0|i52|i0|q i0|i52|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i54|i0|m1 gnd! i0|i54|i0|q i0|i54|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i44|i0|m3 i0|i44|i0|q i0|i44|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i46|i0|m3 i0|i46|i0|q i0|i46|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i52|i0|m3 i0|i52|i0|q i0|i52|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i47|i0|m3 i0|i47|i0|q i0|i47|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i54|i0|m3 i0|i54|i0|q i0|i54|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i44|i0|m11 bl<4> net273 i0|i44|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i46|i0|m11 bl<4> net272 i0|i46|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i52|i0|m11 bl<4> net269 i0|i52|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i54|i0|m11 bl<4> net264 i0|i54|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i45|i3|m10 blb<3> net273 i0|i45|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i47|i3|m10 blb<3> net272 i0|i47|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i53|i3|m10 blb<3> net269 i0|i53|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i55|i3|m10 blb<3> net264 i0|i55|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i45|i3|m1 gnd! i0|i45|i3|q i0|i45|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i53|i0|m3 i0|i53|i0|q i0|i53|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i47|i3|m1 gnd! i0|i47|i3|q i0|i47|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i53|i3|m1 gnd! i0|i53|i3|q i0|i53|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i55|i3|m1 gnd! i0|i55|i3|q i0|i55|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i45|i3|m3 i0|i45|i3|q i0|i45|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i47|i3|m3 i0|i47|i3|q i0|i47|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i53|i3|m3 i0|i53|i3|q i0|i53|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i55|i3|m3 i0|i55|i3|q i0|i55|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i45|i3|m11 bl<3> net273 i0|i45|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i47|i3|m11 bl<3> net272 i0|i47|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i53|i3|m11 bl<3> net269 i0|i53|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i55|i0|m3 i0|i55|i0|q i0|i55|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i55|i3|m11 bl<3> net264 i0|i55|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i45|i2|m10 blb<2> net273 i0|i45|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i47|i2|m10 blb<2> net272 i0|i47|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i53|i2|m10 blb<2> net269 i0|i53|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i55|i2|m10 blb<2> net264 i0|i55|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i45|i2|m1 gnd! i0|i45|i2|q i0|i45|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i47|i2|m1 gnd! i0|i47|i2|q i0|i47|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i53|i2|m1 gnd! i0|i53|i2|q i0|i53|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i55|i2|m1 gnd! i0|i55|i2|q i0|i55|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i45|i2|m3 i0|i45|i2|q i0|i45|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i45|i0|m11 bl<0> net273 i0|i45|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i47|i2|m3 i0|i47|i2|q i0|i47|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i53|i2|m3 i0|i53|i2|q i0|i53|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i55|i2|m3 i0|i55|i2|q i0|i55|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i45|i2|m11 bl<2> net273 i0|i45|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i47|i2|m11 bl<2> net272 i0|i47|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i53|i2|m11 bl<2> net269 i0|i53|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i55|i2|m11 bl<2> net264 i0|i55|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i45|i1|m10 blb<1> net273 i0|i45|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i47|i1|m10 blb<1> net272 i0|i47|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i53|i1|m10 blb<1> net269 i0|i53|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i47|i0|m11 bl<0> net272 i0|i47|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i55|i1|m10 blb<1> net264 i0|i55|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i45|i1|m1 gnd! i0|i45|i1|q i0|i45|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i47|i1|m1 gnd! i0|i47|i1|q i0|i47|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i53|i1|m1 gnd! i0|i53|i1|q i0|i53|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i55|i1|m1 gnd! i0|i55|i1|q i0|i55|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i45|i1|m3 i0|i45|i1|q i0|i45|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i47|i1|m3 i0|i47|i1|q i0|i47|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i53|i1|m3 i0|i53|i1|q i0|i53|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i55|i1|m3 i0|i55|i1|q i0|i55|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i45|i1|m11 bl<1> net273 i0|i45|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i53|i0|m11 bl<0> net269 i0|i53|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i36|i3|m10 blb<7> net277 i0|i36|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i38|i3|m10 blb<7> net276 i0|i38|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i36|i3|m1 gnd! i0|i36|i3|q i0|i36|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i47|i1|m11 bl<1> net272 i0|i47|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i38|i3|m1 gnd! i0|i38|i3|q i0|i38|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i36|i3|m3 i0|i36|i3|q i0|i36|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i38|i3|m3 i0|i38|i3|q i0|i38|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i36|i3|m11 bl<7> net277 i0|i36|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i38|i3|m11 bl<7> net276 i0|i38|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i36|i2|m10 blb<6> net277 i0|i36|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i38|i2|m10 blb<6> net276 i0|i38|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i36|i2|m1 gnd! i0|i36|i2|q i0|i36|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i38|i2|m1 gnd! i0|i38|i2|q i0|i38|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i36|i2|m3 i0|i36|i2|q i0|i36|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i53|i1|m11 bl<1> net269 i0|i53|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i38|i2|m3 i0|i38|i2|q i0|i38|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i36|i2|m11 bl<6> net277 i0|i36|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i38|i2|m11 bl<6> net276 i0|i38|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i36|i1|m10 blb<5> net277 i0|i36|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i38|i1|m10 blb<5> net276 i0|i38|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i36|i1|m1 gnd! i0|i36|i1|q i0|i36|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i38|i1|m1 gnd! i0|i38|i1|q i0|i38|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i36|i1|m3 i0|i36|i1|q i0|i36|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i38|i1|m3 i0|i38|i1|q i0|i38|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i36|i1|m11 bl<5> net277 i0|i36|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i55|i1|m11 bl<1> net264 i0|i55|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i38|i1|m11 bl<5> net276 i0|i38|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i36|i0|m10 blb<4> net277 i0|i36|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i38|i0|m10 blb<4> net276 i0|i38|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i36|i0|m1 gnd! i0|i36|i0|q i0|i36|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i38|i0|m1 gnd! i0|i38|i0|q i0|i38|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i36|i0|m3 i0|i36|i0|q i0|i36|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i38|i0|m3 i0|i38|i0|q i0|i38|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i36|i0|m11 bl<4> net277 i0|i36|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i38|i0|m11 bl<4> net276 i0|i38|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i37|i3|m10 blb<3> net277 i0|i37|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i45|i0|m10 blb<0> net273 i0|i45|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i39|i3|m10 blb<3> net276 i0|i39|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i37|i3|m1 gnd! i0|i37|i3|q i0|i37|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i39|i3|m1 gnd! i0|i39|i3|q i0|i39|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i37|i3|m3 i0|i37|i3|q i0|i37|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i39|i3|m3 i0|i39|i3|q i0|i39|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i37|i3|m11 bl<3> net277 i0|i37|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i39|i3|m11 bl<3> net276 i0|i39|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i37|i2|m10 blb<2> net277 i0|i37|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i39|i2|m10 blb<2> net276 i0|i39|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i37|i2|m1 gnd! i0|i37|i2|q i0|i37|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i47|i0|m10 blb<0> net272 i0|i47|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i39|i2|m1 gnd! i0|i39|i2|q i0|i39|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i37|i2|m3 i0|i37|i2|q i0|i37|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i39|i2|m3 i0|i39|i2|q i0|i39|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i37|i2|m11 bl<2> net277 i0|i37|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i39|i2|m11 bl<2> net276 i0|i39|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i37|i1|m10 blb<1> net277 i0|i37|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i39|i1|m10 blb<1> net276 i0|i39|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i37|i1|m1 gnd! i0|i37|i1|q i0|i37|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i39|i1|m1 gnd! i0|i39|i1|q i0|i39|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i37|i1|m3 i0|i37|i1|q i0|i37|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i53|i0|m10 blb<0> net269 i0|i53|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i39|i1|m3 i0|i39|i1|q i0|i39|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i37|i1|m11 bl<1> net277 i0|i37|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i39|i1|m11 bl<1> net276 i0|i39|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i37|i0|m10 blb<0> net277 i0|i37|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i39|i0|m10 blb<0> net276 i0|i39|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i37|i0|m1 gnd! i0|i37|i0|q i0|i37|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i39|i0|m1 gnd! i0|i39|i0|q i0|i39|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i37|i0|m3 i0|i37|i0|q i0|i37|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i39|i0|m3 i0|i39|i0|q i0|i39|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i37|i0|m11 bl<0> net277 i0|i37|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i55|i0|m10 blb<0> net264 i0|i55|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i39|i0|m11 bl<0> net276 i0|i39|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i44|i3|m10 blb<7> net273 i0|i44|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i46|i3|m10 blb<7> net272 i0|i46|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i52|i3|m10 blb<7> net269 i0|i52|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i54|i3|m10 blb<7> net264 i0|i54|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i44|i3|m1 gnd! i0|i44|i3|q i0|i44|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i46|i3|m1 gnd! i0|i46|i3|q i0|i46|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i52|i3|m1 gnd! i0|i52|i3|q i0|i52|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i54|i3|m1 gnd! i0|i54|i3|q i0|i54|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i44|i3|m3 i0|i44|i3|q i0|i44|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i45|i0|m1 gnd! i0|i45|i0|q i0|i45|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i46|i3|m3 i0|i46|i3|q i0|i46|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i52|i3|m3 i0|i52|i3|q i0|i52|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i54|i3|m3 i0|i54|i3|q i0|i54|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i44|i3|m11 bl<7> net273 i0|i44|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i46|i3|m11 bl<7> net272 i0|i46|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i52|i3|m11 bl<7> net269 i0|i52|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i54|i3|m11 bl<7> net264 i0|i54|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i44|i2|m10 blb<6> net273 i0|i44|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i46|i2|m10 blb<6> net272 i0|i46|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i52|i2|m10 blb<6> net269 i0|i52|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i47|i0|m1 gnd! i0|i47|i0|q i0|i47|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i54|i2|m10 blb<6> net264 i0|i54|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i44|i2|m1 gnd! i0|i44|i2|q i0|i44|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i46|i2|m1 gnd! i0|i46|i2|q i0|i46|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i52|i2|m1 gnd! i0|i52|i2|q i0|i52|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i54|i2|m1 gnd! i0|i54|i2|q i0|i54|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i44|i2|m3 i0|i44|i2|q i0|i44|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i46|i2|m3 i0|i46|i2|q i0|i46|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i52|i2|m3 i0|i52|i2|q i0|i52|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i54|i2|m3 i0|i54|i2|q i0|i54|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i44|i2|m11 bl<6> net273 i0|i44|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i53|i0|m1 gnd! i0|i53|i0|q i0|i53|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i55|i0|m11 bl<0> net264 i0|i55|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i22|i24|m13 gnd! i36|i22|i24|net27 i36|i22|net52 nfet nfin=2 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi36|i22|m4 i36|net269 i36|i22|net52 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i22|i24|m12 ln_x5cbbd88253|x5cbbd882345|17 i36|wen gnd! nfet nfin=2 w=0.021u
+  l=0.015u adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i22|i24|m11 i36|i22|i24|net27 i36|i22|net62 ln_x5cbbd88253|x5cbbd882345|17
+ nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i22|i23|m0 gnd! d<3> i36|i22|net62 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i22|i25|m12 ln_x5cbbd88253|x5cbbd882345|16 d<3> i36|i22|i25|net27 nfet
+ nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi36|i22|i25|m11 gnd! i36|wen ln_x5cbbd88253|x5cbbd882345|16 nfet nfin=2 w=0.021u
+  l=0.015u adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i22|i25|m13 i36|i22|net54 i36|i22|i25|net27 gnd! nfet nfin=2 w=0.021u l=0.015u
+  adeo=2.835e-16 aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i22|m5 i36|net271 i36|i22|net54 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i23|i24|m13 gnd! i36|i23|i24|net27 i36|i23|net52 nfet nfin=2 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi36|i23|m4 i36|net250 i36|i23|net52 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i23|i24|m12 ln_x5cbbd88253|x5cbbd882344|17 i36|wen gnd! nfet nfin=2 w=0.021u
+  l=0.015u adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i23|i24|m11 i36|i23|i24|net27 i36|i23|net62 ln_x5cbbd88253|x5cbbd882344|17
+ nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i23|i23|m0 gnd! d<2> i36|i23|net62 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i23|i25|m12 ln_x5cbbd88253|x5cbbd882344|16 d<2> i36|i23|i25|net27 nfet
+ nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi36|i23|i25|m11 gnd! i36|wen ln_x5cbbd88253|x5cbbd882344|16 nfet nfin=2 w=0.021u
+  l=0.015u adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i23|i25|m13 i36|i23|net54 i36|i23|i25|net27 gnd! nfet nfin=2 w=0.021u l=0.015u
+  adeo=2.835e-16 aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i23|m5 i36|net264 i36|i23|net54 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i24|i24|m13 gnd! i36|i24|i24|net27 i36|i24|net52 nfet nfin=2 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi36|i24|m4 i36|net255 i36|i24|net52 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i24|i24|m12 ln_x5cbbd88253|x5cbbd882343|17 i36|wen gnd! nfet nfin=2 w=0.021u
+  l=0.015u adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i24|i24|m11 i36|i24|i24|net27 i36|i24|net62 ln_x5cbbd88253|x5cbbd882343|17
+ nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i24|i23|m0 gnd! d<1> i36|i24|net62 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i24|i25|m12 ln_x5cbbd88253|x5cbbd882343|16 d<1> i36|i24|i25|net27 nfet
+ nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi36|i24|i25|m11 gnd! i36|wen ln_x5cbbd88253|x5cbbd882343|16 nfet nfin=2 w=0.021u
+  l=0.015u adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i24|i25|m13 i36|i24|net54 i36|i24|i25|net27 gnd! nfet nfin=2 w=0.021u l=0.015u
+  adeo=2.835e-16 aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i24|m5 i36|net263 i36|i24|net54 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i25|i24|m13 gnd! i36|i25|i24|net27 i36|i25|net52 nfet nfin=2 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi36|i25|m4 i36|net254 i36|i25|net52 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i25|i24|m12 ln_x5cbbd88253|x5cbbd882342|17 i36|wen gnd! nfet nfin=2 w=0.021u
+  l=0.015u adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i25|i24|m11 i36|i25|i24|net27 i36|i25|net62 ln_x5cbbd88253|x5cbbd882342|17
+ nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i25|i23|m0 gnd! d<0> i36|i25|net62 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i25|i25|m12 ln_x5cbbd88253|x5cbbd882342|16 d<0> i36|i25|i25|net27 nfet
+ nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi36|i25|i25|m11 gnd! i36|wen ln_x5cbbd88253|x5cbbd882342|16 nfet nfin=2 w=0.021u
+  l=0.015u adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i25|i25|m13 i36|i25|net54 i36|i25|i25|net27 gnd! nfet nfin=2 w=0.021u l=0.015u
+  adeo=2.835e-16 aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i25|m5 i36|net262 i36|i25|net54 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i8|m0 i36|ab<4> a<4> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=2.835e-16
+  pdeo=1.17e-07 pseo=5.85e-08
mi36|i17|m0 i36|wen wenb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=2.835e-16
+  pdeo=1.17e-07 pseo=5.85e-08
mi36|i8|m0@2 gnd! a<4> i36|ab<4> nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i17|m0@2 gnd! wenb i36|wen nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i31|i0|m1 gnd! i0|i31|i0|q i0|i31|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i31|i0|m3 i0|i31|i0|q i0|i31|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i31|i0|m11 bl<0> net280 i0|i31|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi34|i0|i0|m0 i34|i0|net4 net288 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi34|i1|i0|m0 i34|i1|net4 net287 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi34|i2|i0|m0 i34|i2|net4 net286 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi34|i3|i0|m0 i34|i3|net4 net285 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi33|i0|i0|m0 i33|i0|net4 net284 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi33|i1|i0|m0 i33|i1|net4 net283 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi33|i2|i0|m0 i33|i2|net4 net282 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi0|i61|i1|m3 i0|i61|i1|q i0|i61|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi33|i3|i0|m0 i33|i3|net4 net281 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi32|i0|i0|m0 i32|i0|net4 net268 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi32|i1|i0|m0 i32|i1|net4 net267 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi32|i2|i0|m0 i32|i2|net4 net266 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi32|i3|i0|m0 i32|i3|net4 net265 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi34|i0|i0|m0@2 gnd! net288 i34|i0|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi34|i1|i0|m0@2 gnd! net287 i34|i1|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi34|i2|i0|m0@2 gnd! net286 i34|i2|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi34|i3|i0|m0@2 gnd! net285 i34|i3|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi33|i0|i0|m0@2 gnd! net284 i33|i0|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i28|m1 i36|net254 i36|ab<4> bl<0> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi33|i1|i0|m0@2 gnd! net283 i33|i1|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi33|i2|i0|m0@2 gnd! net282 i33|i2|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi33|i3|i0|m0@2 gnd! net281 i33|i3|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi32|i0|i0|m0@2 gnd! net268 i32|i0|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi32|i1|i0|m0@2 gnd! net267 i32|i1|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi32|i2|i0|m0@2 gnd! net266 i32|i2|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi32|i3|i0|m0@2 gnd! net265 i32|i3|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi34|i0|i1|m0 net276 i34|i0|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi34|i1|i1|m0 net275 i34|i1|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi34|i2|i1|m0 net274 i34|i2|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi0|i61|i1|m11 bl<1> net261 i0|i61|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi34|i3|i1|m0 net273 i34|i3|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi33|i0|i1|m0 net272 i33|i0|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi33|i1|i1|m0 net271 i33|i1|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi33|i2|i1|m0 net270 i33|i2|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi33|i3|i1|m0 net269 i33|i3|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi32|i0|i1|m0 net264 i32|i0|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi32|i1|i1|m0 net263 i32|i1|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi32|i2|i1|m0 net262 i32|i2|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi32|i3|i1|m0 net261 i32|i3|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi34|i0|i1|m0@2 gnd! i34|i0|net4 net276 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i61|i0|m10 blb<0> net261 i0|i61|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi34|i1|i1|m0@2 gnd! i34|i1|net4 net275 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi34|i2|i1|m0@2 gnd! i34|i2|net4 net274 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi34|i3|i1|m0@2 gnd! i34|i3|net4 net273 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi33|i0|i1|m0@2 gnd! i33|i0|net4 net272 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi33|i1|i1|m0@2 gnd! i33|i1|net4 net271 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi33|i2|i1|m0@2 gnd! i33|i2|net4 net270 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi33|i3|i1|m0@2 gnd! i33|i3|net4 net269 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi32|i0|i1|m0@2 gnd! i32|i0|net4 net264 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi32|i1|i1|m0@2 gnd! i32|i1|net4 net263 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi32|i2|i1|m0@2 gnd! i32|i2|net4 net262 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i32|m0 i36|net262 a<4> blb<4> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi32|i3|i1|m0@2 gnd! i32|i3|net4 net261 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i60|i3|m10 blb<7> net261 i0|i60|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i26|m0 i36|net269 a<4> bl<7> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i3|m1 gnd! i0|i60|i3|q i0|i60|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i3|m3 i0|i60|i3|q i0|i60|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i26|m1 i36|net269 i36|ab<4> bl<3> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i3|m11 bl<7> net261 i0|i60|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i60|i2|m10 blb<6> net261 i0|i60|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i29|m0 i36|net271 a<4> blb<7> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i2|m1 gnd! i0|i60|i2|q i0|i60|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i61|i0|m1 gnd! i0|i61|i0|q i0|i61|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i2|m3 i0|i60|i2|q i0|i60|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i29|m1 i36|net271 i36|ab<4> blb<3> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i2|m11 bl<6> net261 i0|i60|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i60|i1|m10 blb<5> net261 i0|i60|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i9|m0 i36|net250 a<4> bl<6> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i1|m1 gnd! i0|i60|i1|q i0|i60|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i1|m3 i0|i60|i1|q i0|i60|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i9|m1 i36|net250 i36|ab<4> bl<2> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i1|m11 bl<5> net261 i0|i60|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i60|i0|m10 blb<4> net261 i0|i60|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i61|i0|m3 i0|i61|i0|q i0|i61|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i30|m0 i36|net264 a<4> blb<6> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i0|m1 gnd! i0|i60|i0|q i0|i60|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i0|m3 i0|i60|i0|q i0|i60|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i30|m1 i36|net264 i36|ab<4> blb<2> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i60|i0|m11 bl<4> net261 i0|i60|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i61|i3|m10 blb<3> net261 i0|i61|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi36|i27|m0 i36|net255 a<4> bl<5> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i61|i3|m1 gnd! i0|i61|i3|q i0|i61|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i61|i3|m3 i0|i61|i3|q i0|i61|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i27|m1 i36|net255 i36|ab<4> bl<1> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i32|m1 i36|net262 i36|ab<4> blb<0> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i61|i3|m11 bl<3> net261 i0|i61|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i61|i2|m10 blb<2> net261 i0|i61|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi11|m188 net291 i11|net697 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=2.835e-16 pdeo=5.85e-08 pseo=5.85e-08
mi36|i31|m0 i36|net263 a<4> blb<5> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi11|m117 net291 a<1> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m104 net291 a<2> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m93 net291 a<3> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m131 net292 a<0> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m116 net292 a<1> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m103 net292 a<2> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi11|m94 net292 a<3> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=2.835e-16
+  pdeo=5.85e-08 pseo=5.85e-08
mi35|i0|i0|m0 i35|i0|net4 net292 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi35|i1|i0|m0 i35|i1|net4 net291 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi35|i2|i0|m0 i35|i2|net4 net290 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi0|i61|i2|m1 gnd! i0|i61|i2|q i0|i61|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi35|i3|i0|m0 i35|i3|net4 net289 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi35|i0|i0|m0@2 gnd! net292 i35|i0|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi35|i1|i0|m0@2 gnd! net291 i35|i1|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi35|i2|i0|m0@2 gnd! net290 i35|i2|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi35|i3|i0|m0@2 gnd! net289 i35|i3|net4 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi39|i30|m0 i39|ab<4> a<4> gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi35|i0|i1|m0 net280 i35|i0|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi35|i1|i1|m0 net279 i35|i1|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi35|i2|i1|m0 net278 i35|i2|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi35|i3|i1|m0 net277 i35|i3|net4 gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi0|i61|i2|m3 i0|i61|i2|q i0|i61|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi39|i30|m0@2 gnd! a<4> i39|ab<4> nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+ aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi35|i0|i1|m0@2 gnd! i35|i0|net4 net280 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi35|i1|i1|m0@2 gnd! i35|i1|net4 net279 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi35|i2|i1|m0@2 gnd! i35|i2|net4 net278 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi35|i3|i1|m0@2 gnd! i35|i3|net4 net277 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i30|i3|m10 blb<7> net280 i0|i30|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i30|i3|m1 gnd! i0|i30|i3|q i0|i30|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i30|i3|m3 i0|i30|i3|q i0|i30|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i30|i3|m11 bl<7> net280 i0|i30|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi39|i22|m3 ln_156 wenb bl<7> nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=2.835e-16
+  pdeo=1.17e-07 pseo=5.85e-08
mi36|i31|m1 i36|net263 i36|ab<4> blb<1> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi39|i22|m0 net229 a<4> ln_156 nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi39|i22|m2 ln_157 i39|ab<4> net229 nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i30|i2|m10 blb<6> net280 i0|i30|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi39|i22|m1 bl<3> wenb ln_157 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=5.67e-16
+  pdeo=5.85e-08 pseo=1.17e-07
mi0|i30|i2|m1 gnd! i0|i30|i2|q i0|i30|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i30|i2|m3 i0|i30|i2|q i0|i30|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i30|i2|m11 bl<6> net280 i0|i30|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i30|i1|m10 blb<5> net280 i0|i30|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i30|i1|m1 gnd! i0|i30|i1|q i0|i30|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i30|i1|m3 i0|i30|i1|q i0|i30|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i61|i2|m11 bl<2> net261 i0|i61|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi39|i23|m3 ln_154 wenb bl<6> nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=2.835e-16
+  pdeo=1.17e-07 pseo=5.85e-08
mi0|i30|i1|m11 bl<5> net280 i0|i30|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi39|i23|m0 net227 a<4> ln_154 nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi39|i23|m2 ln_155 i39|ab<4> net227 nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi39|i23|m1 bl<2> wenb ln_155 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=5.67e-16
+  pdeo=5.85e-08 pseo=1.17e-07
mi0|i30|i0|m10 blb<4> net280 i0|i30|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i30|i0|m1 gnd! i0|i30|i0|q i0|i30|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i30|i0|m3 i0|i30|i0|q i0|i30|i0|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i30|i0|m11 bl<4> net280 i0|i30|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i31|i3|m10 blb<3> net280 i0|i31|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i61|i1|m10 blb<1> net261 i0|i61|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i31|i3|m1 gnd! i0|i31|i3|q i0|i31|i3|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i31|i3|m3 i0|i31|i3|q i0|i31|i3|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi39|i24|m3 ln_152 wenb bl<5> nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=2.835e-16
+  pdeo=1.17e-07 pseo=5.85e-08
mi0|i31|i3|m11 bl<3> net280 i0|i31|i3|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi39|i24|m0 net225 a<4> ln_152 nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi39|i24|m2 ln_153 i39|ab<4> net225 nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi39|i24|m1 bl<1> wenb ln_153 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=5.67e-16
+  pdeo=5.85e-08 pseo=1.17e-07
mi0|i31|i2|m10 blb<2> net280 i0|i31|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i31|i2|m1 gnd! i0|i31|i2|q i0|i31|i2|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i31|i2|m3 i0|i31|i2|q i0|i31|i2|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i28|m0 i36|net254 a<4> bl<4> nfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i31|i2|m11 bl<2> net280 i0|i31|i2|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i31|i1|m10 blb<1> net280 i0|i31|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i31|i1|m1 gnd! i0|i31|i1|q i0|i31|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i31|i1|m3 i0|i31|i1|q i0|i31|i1|qb gnd! nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi39|i25|m3 ln_150 wenb bl<4> nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=2.835e-16
+  pdeo=1.17e-07 pseo=5.85e-08
mi0|i31|i1|m11 bl<1> net280 i0|i31|i1|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi39|i25|m0 net355 a<4> ln_150 nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi39|i25|m2 ln_151 i39|ab<4> net355 nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi39|i25|m1 bl<0> wenb ln_151 nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16 aseo=5.67e-16
+  pdeo=5.85e-08 pseo=1.17e-07
mi0|i31|i0|m10 blb<0> net280 i0|i31|i0|qb nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi0|i61|i1|m1 gnd! i0|i61|i1|q i0|i61|i1|qb nfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi0|i61|i0|m11 bl<0> net261 i0|i61|i0|q nfet nfin=2 w=0.021u l=0.015u adeo=2.835e-16
+  aseo=5.67e-16 pdeo=5.85e-08 pseo=1.17e-07
mi11|m12 net268 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m14 net266 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m8 net284 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m10 net282 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m4 net288 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m6 net286 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m0 net292 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m2 net290 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m13 net267 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m15 net265 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m9 net283 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m11 net281 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m5 net287 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m7 net285 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m1 net291 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi11|m3 net289 clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=5.67e-16
+  pdeo=1.17e-07 pseo=1.17e-07
mi0|i61|i2|m4 i0|i61|i2|q i0|i61|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i59|i1|m2 i0|i59|i1|qb i0|i59|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i61|i1|m2 i0|i61|i1|qb i0|i61|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i59|i1|m4 i0|i59|i1|q i0|i59|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i61|i1|m4 i0|i61|i1|q i0|i61|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i59|i0|m2 i0|i59|i0|qb i0|i59|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i61|i0|m2 i0|i61|i0|qb i0|i61|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i59|i0|m4 i0|i59|i0|q i0|i59|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i59|i3|m2 i0|i59|i3|qb i0|i59|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i61|i3|m2 i0|i61|i3|qb i0|i61|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i59|i3|m4 i0|i59|i3|q i0|i59|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i61|i3|m4 i0|i61|i3|q i0|i61|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i59|i2|m2 i0|i59|i2|qb i0|i59|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i61|i2|m2 i0|i61|i2|qb i0|i61|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i59|i2|m4 i0|i59|i2|q i0|i59|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i61|i0|m4 i0|i61|i0|q i0|i61|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i57|i2|m4 i0|i57|i2|q i0|i57|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i55|i1|m2 i0|i55|i1|qb i0|i55|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i57|i1|m2 i0|i57|i1|qb i0|i57|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i55|i1|m4 i0|i55|i1|q i0|i55|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i57|i1|m4 i0|i57|i1|q i0|i57|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i55|i0|m2 i0|i55|i0|qb i0|i55|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i57|i0|m2 i0|i57|i0|qb i0|i57|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i55|i0|m4 i0|i55|i0|q i0|i55|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i55|i3|m2 i0|i55|i3|qb i0|i55|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i57|i3|m2 i0|i57|i3|qb i0|i57|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i55|i3|m4 i0|i55|i3|q i0|i55|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i57|i3|m4 i0|i57|i3|q i0|i57|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i55|i2|m2 i0|i55|i2|qb i0|i55|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i57|i2|m2 i0|i57|i2|qb i0|i57|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i55|i2|m4 i0|i55|i2|q i0|i55|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i57|i0|m4 i0|i57|i0|q i0|i57|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i53|i2|m4 i0|i53|i2|q i0|i53|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i51|i1|m2 i0|i51|i1|qb i0|i51|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i53|i1|m2 i0|i53|i1|qb i0|i53|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i51|i1|m4 i0|i51|i1|q i0|i51|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i53|i1|m4 i0|i53|i1|q i0|i53|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i51|i0|m2 i0|i51|i0|qb i0|i51|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i53|i0|m2 i0|i53|i0|qb i0|i53|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i51|i0|m4 i0|i51|i0|q i0|i51|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i51|i3|m2 i0|i51|i3|qb i0|i51|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i53|i3|m2 i0|i53|i3|qb i0|i53|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i51|i3|m4 i0|i51|i3|q i0|i51|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i53|i3|m4 i0|i53|i3|q i0|i53|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i51|i2|m2 i0|i51|i2|qb i0|i51|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i53|i2|m2 i0|i53|i2|qb i0|i53|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i51|i2|m4 i0|i51|i2|q i0|i51|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i53|i0|m4 i0|i53|i0|q i0|i53|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i49|i2|m4 i0|i49|i2|q i0|i49|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i47|i1|m2 i0|i47|i1|qb i0|i47|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i49|i1|m2 i0|i49|i1|qb i0|i49|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i47|i1|m4 i0|i47|i1|q i0|i47|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i49|i1|m4 i0|i49|i1|q i0|i49|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i47|i0|m2 i0|i47|i0|qb i0|i47|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i49|i0|m2 i0|i49|i0|qb i0|i49|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i47|i0|m4 i0|i47|i0|q i0|i47|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i47|i3|m2 i0|i47|i3|qb i0|i47|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i49|i3|m2 i0|i49|i3|qb i0|i49|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i47|i3|m4 i0|i47|i3|q i0|i47|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i49|i3|m4 i0|i49|i3|q i0|i49|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i47|i2|m2 i0|i47|i2|qb i0|i47|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i49|i2|m2 i0|i49|i2|qb i0|i49|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i47|i2|m4 i0|i47|i2|q i0|i47|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i49|i0|m4 i0|i49|i0|q i0|i49|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i45|i2|m4 i0|i45|i2|q i0|i45|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i43|i1|m2 i0|i43|i1|qb i0|i43|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i45|i1|m2 i0|i45|i1|qb i0|i45|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i43|i1|m4 i0|i43|i1|q i0|i43|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i45|i1|m4 i0|i45|i1|q i0|i45|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i43|i0|m2 i0|i43|i0|qb i0|i43|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i45|i0|m2 i0|i45|i0|qb i0|i45|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i43|i0|m4 i0|i43|i0|q i0|i43|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i43|i3|m2 i0|i43|i3|qb i0|i43|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i45|i3|m2 i0|i45|i3|qb i0|i45|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i43|i3|m4 i0|i43|i3|q i0|i43|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i45|i3|m4 i0|i45|i3|q i0|i45|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i43|i2|m2 i0|i43|i2|qb i0|i43|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i45|i2|m2 i0|i45|i2|qb i0|i45|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i43|i2|m4 i0|i43|i2|q i0|i43|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i45|i0|m4 i0|i45|i0|q i0|i45|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i41|i2|m4 i0|i41|i2|q i0|i41|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i39|i1|m2 i0|i39|i1|qb i0|i39|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i41|i1|m2 i0|i41|i1|qb i0|i41|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i39|i1|m4 i0|i39|i1|q i0|i39|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i41|i1|m4 i0|i41|i1|q i0|i41|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i39|i0|m2 i0|i39|i0|qb i0|i39|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i41|i0|m2 i0|i41|i0|qb i0|i41|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i39|i0|m4 i0|i39|i0|q i0|i39|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i39|i3|m2 i0|i39|i3|qb i0|i39|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i41|i3|m2 i0|i41|i3|qb i0|i41|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i39|i3|m4 i0|i39|i3|q i0|i39|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i41|i3|m4 i0|i41|i3|q i0|i41|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i39|i2|m2 i0|i39|i2|qb i0|i39|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i41|i2|m2 i0|i41|i2|qb i0|i41|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i39|i2|m4 i0|i39|i2|q i0|i39|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i41|i0|m4 i0|i41|i0|q i0|i41|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i37|i2|m4 i0|i37|i2|q i0|i37|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i35|i1|m2 i0|i35|i1|qb i0|i35|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i37|i1|m2 i0|i37|i1|qb i0|i37|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i35|i1|m4 i0|i35|i1|q i0|i35|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i37|i1|m4 i0|i37|i1|q i0|i37|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i35|i0|m2 i0|i35|i0|qb i0|i35|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i37|i0|m2 i0|i37|i0|qb i0|i37|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i35|i0|m4 i0|i35|i0|q i0|i35|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i35|i3|m2 i0|i35|i3|qb i0|i35|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i37|i3|m2 i0|i37|i3|qb i0|i37|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i35|i3|m4 i0|i35|i3|q i0|i35|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i37|i3|m4 i0|i37|i3|q i0|i37|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i35|i2|m2 i0|i35|i2|qb i0|i35|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i37|i2|m2 i0|i37|i2|qb i0|i37|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i35|i2|m4 i0|i35|i2|q i0|i35|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i37|i0|m4 i0|i37|i0|q i0|i37|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i33|i2|m4 i0|i33|i2|q i0|i33|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i31|i1|m2 i0|i31|i1|qb i0|i31|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i33|i1|m2 i0|i33|i1|qb i0|i33|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i31|i1|m4 i0|i31|i1|q i0|i31|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i33|i1|m4 i0|i33|i1|q i0|i33|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i31|i0|m2 i0|i31|i0|qb i0|i31|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i33|i0|m2 i0|i33|i0|qb i0|i33|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i31|i0|m4 i0|i31|i0|q i0|i31|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i31|i3|m2 i0|i31|i3|qb i0|i31|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i33|i3|m2 i0|i33|i3|qb i0|i33|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i31|i3|m4 i0|i31|i3|q i0|i31|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i33|i3|m4 i0|i33|i3|q i0|i33|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i31|i2|m2 i0|i31|i2|qb i0|i31|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i33|i2|m2 i0|i33|i2|qb i0|i33|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i31|i2|m4 i0|i31|i2|q i0|i31|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i33|i0|m4 i0|i33|i0|q i0|i33|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i60|i2|m4 i0|i60|i2|q i0|i60|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i58|i1|m2 i0|i58|i1|qb i0|i58|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i60|i1|m2 i0|i60|i1|qb i0|i60|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i58|i1|m4 i0|i58|i1|q i0|i58|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i60|i1|m4 i0|i60|i1|q i0|i60|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i58|i0|m2 i0|i58|i0|qb i0|i58|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i60|i0|m2 i0|i60|i0|qb i0|i60|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i58|i0|m4 i0|i58|i0|q i0|i58|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i58|i3|m2 i0|i58|i3|qb i0|i58|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i60|i3|m2 i0|i60|i3|qb i0|i60|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i58|i3|m4 i0|i58|i3|q i0|i58|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i60|i3|m4 i0|i60|i3|q i0|i60|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i58|i2|m2 i0|i58|i2|qb i0|i58|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i60|i2|m2 i0|i60|i2|qb i0|i60|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i58|i2|m4 i0|i58|i2|q i0|i58|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i60|i0|m4 i0|i60|i0|q i0|i60|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i56|i2|m4 i0|i56|i2|q i0|i56|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i54|i1|m2 i0|i54|i1|qb i0|i54|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i56|i1|m2 i0|i56|i1|qb i0|i56|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i54|i1|m4 i0|i54|i1|q i0|i54|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i56|i1|m4 i0|i56|i1|q i0|i56|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i54|i0|m2 i0|i54|i0|qb i0|i54|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i56|i0|m2 i0|i56|i0|qb i0|i56|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i54|i0|m4 i0|i54|i0|q i0|i54|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i54|i3|m2 i0|i54|i3|qb i0|i54|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i56|i3|m2 i0|i56|i3|qb i0|i56|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i54|i3|m4 i0|i54|i3|q i0|i54|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i56|i3|m4 i0|i56|i3|q i0|i56|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i54|i2|m2 i0|i54|i2|qb i0|i54|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i56|i2|m2 i0|i56|i2|qb i0|i56|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i54|i2|m4 i0|i54|i2|q i0|i54|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i56|i0|m4 i0|i56|i0|q i0|i56|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i52|i2|m4 i0|i52|i2|q i0|i52|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i50|i1|m2 i0|i50|i1|qb i0|i50|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i52|i1|m2 i0|i52|i1|qb i0|i52|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i50|i1|m4 i0|i50|i1|q i0|i50|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i52|i1|m4 i0|i52|i1|q i0|i52|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i50|i0|m2 i0|i50|i0|qb i0|i50|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i52|i0|m2 i0|i52|i0|qb i0|i52|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i50|i0|m4 i0|i50|i0|q i0|i50|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i50|i3|m2 i0|i50|i3|qb i0|i50|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i52|i3|m2 i0|i52|i3|qb i0|i52|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i50|i3|m4 i0|i50|i3|q i0|i50|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i52|i3|m4 i0|i52|i3|q i0|i52|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i50|i2|m2 i0|i50|i2|qb i0|i50|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i52|i2|m2 i0|i52|i2|qb i0|i52|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i50|i2|m4 i0|i50|i2|q i0|i50|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i52|i0|m4 i0|i52|i0|q i0|i52|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i48|i2|m4 i0|i48|i2|q i0|i48|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i46|i1|m2 i0|i46|i1|qb i0|i46|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i48|i1|m2 i0|i48|i1|qb i0|i48|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i46|i1|m4 i0|i46|i1|q i0|i46|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i48|i1|m4 i0|i48|i1|q i0|i48|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i46|i0|m2 i0|i46|i0|qb i0|i46|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i48|i0|m2 i0|i48|i0|qb i0|i48|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i46|i0|m4 i0|i46|i0|q i0|i46|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i46|i3|m2 i0|i46|i3|qb i0|i46|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i48|i3|m2 i0|i48|i3|qb i0|i48|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i46|i3|m4 i0|i46|i3|q i0|i46|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i48|i3|m4 i0|i48|i3|q i0|i48|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i46|i2|m2 i0|i46|i2|qb i0|i46|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i48|i2|m2 i0|i48|i2|qb i0|i48|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i46|i2|m4 i0|i46|i2|q i0|i46|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i48|i0|m4 i0|i48|i0|q i0|i48|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i44|i2|m4 i0|i44|i2|q i0|i44|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i42|i1|m2 i0|i42|i1|qb i0|i42|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i44|i1|m2 i0|i44|i1|qb i0|i44|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i42|i1|m4 i0|i42|i1|q i0|i42|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i44|i1|m4 i0|i44|i1|q i0|i44|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i42|i0|m2 i0|i42|i0|qb i0|i42|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i44|i0|m2 i0|i44|i0|qb i0|i44|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i42|i0|m4 i0|i42|i0|q i0|i42|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i42|i3|m2 i0|i42|i3|qb i0|i42|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i44|i3|m2 i0|i44|i3|qb i0|i44|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i42|i3|m4 i0|i42|i3|q i0|i42|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i44|i3|m4 i0|i44|i3|q i0|i44|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i42|i2|m2 i0|i42|i2|qb i0|i42|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i44|i2|m2 i0|i44|i2|qb i0|i44|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i42|i2|m4 i0|i42|i2|q i0|i42|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i44|i0|m4 i0|i44|i0|q i0|i44|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i40|i2|m4 i0|i40|i2|q i0|i40|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i38|i1|m2 i0|i38|i1|qb i0|i38|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i40|i1|m2 i0|i40|i1|qb i0|i40|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i38|i1|m4 i0|i38|i1|q i0|i38|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i40|i1|m4 i0|i40|i1|q i0|i40|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i38|i0|m2 i0|i38|i0|qb i0|i38|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i40|i0|m2 i0|i40|i0|qb i0|i40|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i38|i0|m4 i0|i38|i0|q i0|i38|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i38|i3|m2 i0|i38|i3|qb i0|i38|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i40|i3|m2 i0|i40|i3|qb i0|i40|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i38|i3|m4 i0|i38|i3|q i0|i38|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i40|i3|m4 i0|i40|i3|q i0|i40|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i38|i2|m2 i0|i38|i2|qb i0|i38|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i40|i2|m2 i0|i40|i2|qb i0|i40|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i38|i2|m4 i0|i38|i2|q i0|i38|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i40|i0|m4 i0|i40|i0|q i0|i40|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i36|i2|m4 i0|i36|i2|q i0|i36|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i34|i1|m2 i0|i34|i1|qb i0|i34|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i36|i1|m2 i0|i36|i1|qb i0|i36|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i34|i1|m4 i0|i34|i1|q i0|i34|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i36|i1|m4 i0|i36|i1|q i0|i36|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i34|i0|m2 i0|i34|i0|qb i0|i34|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i36|i0|m2 i0|i36|i0|qb i0|i36|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i34|i0|m4 i0|i34|i0|q i0|i34|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i34|i3|m2 i0|i34|i3|qb i0|i34|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i36|i3|m2 i0|i36|i3|qb i0|i36|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i34|i3|m4 i0|i34|i3|q i0|i34|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i36|i3|m4 i0|i36|i3|q i0|i36|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i34|i2|m2 i0|i34|i2|qb i0|i34|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i36|i2|m2 i0|i36|i2|qb i0|i36|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i34|i2|m4 i0|i34|i2|q i0|i34|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i36|i0|m4 i0|i36|i0|q i0|i36|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i32|i2|m4 i0|i32|i2|q i0|i32|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i30|i1|m2 i0|i30|i1|qb i0|i30|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i32|i1|m2 i0|i32|i1|qb i0|i32|i1|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i30|i1|m4 i0|i30|i1|q i0|i30|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i32|i1|m4 i0|i32|i1|q i0|i32|i1|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i30|i0|m2 i0|i30|i0|qb i0|i30|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i32|i0|m2 i0|i32|i0|qb i0|i32|i0|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i30|i0|m4 i0|i30|i0|q i0|i30|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i30|i3|m2 i0|i30|i3|qb i0|i30|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i32|i3|m2 i0|i32|i3|qb i0|i32|i3|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i30|i3|m4 i0|i30|i3|q i0|i30|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i32|i3|m4 i0|i32|i3|q i0|i32|i3|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i30|i2|m2 i0|i30|i2|qb i0|i30|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i32|i2|m2 i0|i32|i2|qb i0|i32|i2|q vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i30|i2|m4 i0|i30|i2|q i0|i30|i2|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi0|i32|i0|m4 i0|i32|i0|q i0|i32|i0|qb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi36|i22|i24|m14 i36|i22|i24|net27 i36|i22|net62 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=1.134e-15 aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi36|i22|i24|m15 vdd! i36|wen i36|i22|i24|net27 pfet nfin=4 w=0.021u l=0.015u
+ adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
mi36|i22|i24|m16 i36|i22|net52 i36|i22|i24|net27 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi36|i22|i25|m14 i36|i22|i25|net27 d<3> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi36|i22|i25|m15 vdd! i36|wen i36|i22|i25|net27 pfet nfin=4 w=0.021u l=0.015u
+ adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
mi36|i22|i25|m16 i36|i22|net54 i36|i22|i25|net27 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi36|i22|i23|m1 i36|i22|net62 d<3> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i23|i24|m14 i36|i23|i24|net27 i36|i23|net62 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=1.134e-15 aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi36|i23|i24|m15 vdd! i36|wen i36|i23|i24|net27 pfet nfin=4 w=0.021u l=0.015u
+ adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
mi36|i23|i24|m16 i36|i23|net52 i36|i23|i24|net27 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi36|i23|i25|m15 i36|i23|i25|net27 d<2> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi36|i23|i25|m14 vdd! i36|wen i36|i23|i25|net27 pfet nfin=4 w=0.021u l=0.015u
+ adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
mi36|i23|i25|m16 i36|i23|net54 i36|i23|i25|net27 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi36|i23|i23|m1 i36|i23|net62 d<2> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i24|i24|m14 i36|i24|i24|net27 i36|i24|net62 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=1.134e-15 aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi36|i24|i24|m15 vdd! i36|wen i36|i24|i24|net27 pfet nfin=4 w=0.021u l=0.015u
+ adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
mi36|i24|i24|m16 i36|i24|net52 i36|i24|i24|net27 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi36|i24|i25|m15 i36|i24|i25|net27 d<1> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi36|i24|i25|m14 vdd! i36|wen i36|i24|i25|net27 pfet nfin=4 w=0.021u l=0.015u
+ adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
mi36|i24|i25|m16 i36|i24|net54 i36|i24|i25|net27 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi36|i24|i23|m1 i36|i24|net62 d<1> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i25|i24|m14 i36|i25|i24|net27 i36|i25|net62 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=1.134e-15 aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi36|i25|i24|m15 vdd! i36|wen i36|i25|i24|net27 pfet nfin=4 w=0.021u l=0.015u
+ adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
mi36|i25|i24|m16 i36|i25|net52 i36|i25|i24|net27 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi36|i25|i25|m15 i36|i25|i25|net27 d<0> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi36|i25|i25|m14 vdd! i36|wen i36|i25|i25|net27 pfet nfin=4 w=0.021u l=0.015u
+ adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
mi36|i25|i25|m16 i36|i25|net54 i36|i25|i25|net27 vdd! pfet nfin=4 w=0.021u l=0.015u
+  adeo=5.67e-16 aseo=1.134e-15 pdeo=1.17e-07 pseo=2.34e-07
mi36|i25|i23|m1 i36|i25|net62 d<0> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16
+  aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
mi36|i8|m1 i36|ab<4> a<4> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+ aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi36|i17|m1 i36|wen wenb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi36|i8|m1@2 i36|ab<4> a<4> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+ aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi36|i17|m1@2 i36|wen wenb vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+ aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi6|i1|m2 bl<1> clk blb<1> pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i0|m0@2 blb<0> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i1|m2@2 bl<1> clk blb<1> pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i1|m1 bl<1> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i0|m2 bl<0> clk blb<0> pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i7|m0 blb<7> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i7|m0@2 blb<7> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i6|m0 blb<6> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i7|m2 bl<7> clk blb<7> pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i6|m0@2 blb<6> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i7|m2@2 bl<7> clk blb<7> pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i7|m1 bl<7> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i6|m2 bl<6> clk blb<6> pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i7|m1@2 bl<7> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i1|m1@2 bl<1> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i6|m2@2 bl<6> clk blb<6> pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i6|m1 bl<6> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i6|m1@2 bl<6> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i5|m0 blb<5> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i5|m0@2 blb<5> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i4|m0 blb<4> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i5|m2 bl<5> clk blb<5> pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i4|m0@2 blb<4> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i5|m2@2 bl<5> clk blb<5> pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i5|m1 bl<5> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i0|m2@2 bl<0> clk blb<0> pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i4|m2 bl<4> clk blb<4> pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i5|m1@2 bl<5> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i4|m2@2 bl<4> clk blb<4> pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i4|m1 bl<4> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i4|m1@2 bl<4> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i3|m0 blb<3> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i3|m0@2 blb<3> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i2|m0 blb<2> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i3|m2 bl<3> clk blb<3> pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i2|m0@2 blb<2> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i0|m1 bl<0> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i3|m2@2 bl<3> clk blb<3> pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i3|m1 bl<3> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i2|m2 bl<2> clk blb<2> pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i3|m1@2 bl<3> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i2|m2@2 bl<2> clk blb<2> pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i2|m1 bl<2> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=1.134e-15
+  pdeo=2.34e-07 pseo=2.34e-07
mi6|i2|m1@2 bl<2> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi6|i1|m0 blb<1> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i1|m0@2 blb<1> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i0|m0 blb<0> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15 aseo=5.67e-16
+  pdeo=2.34e-07 pseo=1.17e-07
mi6|i0|m1@2 bl<0> clk vdd! pfet nfin=4 w=0.021u l=0.015u adeo=5.67e-16 aseo=1.134e-15
+  pdeo=1.17e-07 pseo=2.34e-07
mi11|i232|m1 i11|net697 a<0> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+ aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi11|i232|m1@2 i11|net697 a<0> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi11|i233|m1 i11|net698 a<1> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+ aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi11|i233|m1@2 i11|net698 a<1> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi11|i234|m1 i11|net699 a<2> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+ aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi11|i234|m1@2 i11|net699 a<2> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi11|i235|m1 i11|net700 a<3> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+ aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi11|i235|m1@2 i11|net700 a<3> vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i0|i0|m1 i35|i0|net4 net292 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i1|i0|m1 i35|i1|net4 net291 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i2|i0|m1 i35|i2|net4 net290 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i3|i0|m1 i35|i3|net4 net289 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i0|i0|m1 i34|i0|net4 net288 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i1|i0|m1 i34|i1|net4 net287 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i2|i0|m1 i34|i2|net4 net286 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i3|i0|m1 i34|i3|net4 net285 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i0|i0|m1 i33|i0|net4 net284 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i1|i0|m1 i33|i1|net4 net283 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i2|i0|m1 i33|i2|net4 net282 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i3|i0|m1 i33|i3|net4 net281 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i0|i0|m1 i32|i0|net4 net268 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i1|i0|m1 i32|i1|net4 net267 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i2|i0|m1 i32|i2|net4 net266 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i3|i0|m1 i32|i3|net4 net265 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i0|i0|m1@2 i35|i0|net4 net292 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i1|i0|m1@2 i35|i1|net4 net291 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i2|i0|m1@2 i35|i2|net4 net290 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i3|i0|m1@2 i35|i3|net4 net289 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i0|i0|m1@2 i34|i0|net4 net288 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i1|i0|m1@2 i34|i1|net4 net287 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i2|i0|m1@2 i34|i2|net4 net286 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i3|i0|m1@2 i34|i3|net4 net285 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i0|i0|m1@2 i33|i0|net4 net284 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i1|i0|m1@2 i33|i1|net4 net283 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i2|i0|m1@2 i33|i2|net4 net282 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i3|i0|m1@2 i33|i3|net4 net281 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i0|i0|m1@2 i32|i0|net4 net268 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i1|i0|m1@2 i32|i1|net4 net267 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i2|i0|m1@2 i32|i2|net4 net266 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i3|i0|m1@2 i32|i3|net4 net265 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi39|i30|m1 i39|ab<4> a<4> vdd! pfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi35|i0|i1|m1 net280 i35|i0|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i1|i1|m1 net279 i35|i1|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i2|i1|m1 net278 i35|i2|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i3|i1|m1 net277 i35|i3|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i0|i1|m1 net276 i34|i0|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i1|i1|m1 net275 i34|i1|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i2|i1|m1 net274 i34|i2|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i3|i1|m1 net273 i34|i3|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i0|i1|m1 net272 i33|i0|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i1|i1|m1 net271 i33|i1|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i2|i1|m1 net270 i33|i2|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i3|i1|m1 net269 i33|i3|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i0|i1|m1 net264 i32|i0|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i1|i1|m1 net263 i32|i1|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i2|i1|m1 net262 i32|i2|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i3|i1|m1 net261 i32|i3|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi39|i30|m1@2 i39|ab<4> a<4> vdd! pfet nfin=2 w=0.021u l=0.015u adeo=5.67e-16
+ aseo=2.835e-16 pdeo=1.17e-07 pseo=5.85e-08
mi35|i0|i1|m1@2 net280 i35|i0|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i1|i1|m1@2 net279 i35|i1|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i2|i1|m1@2 net278 i35|i2|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi35|i3|i1|m1@2 net277 i35|i3|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i0|i1|m1@2 net276 i34|i0|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i1|i1|m1@2 net275 i34|i1|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i2|i1|m1@2 net274 i34|i2|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi34|i3|i1|m1@2 net273 i34|i3|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i0|i1|m1@2 net272 i33|i0|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i1|i1|m1@2 net271 i33|i1|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i2|i1|m1@2 net270 i33|i2|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi33|i3|i1|m1@2 net269 i33|i3|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i0|i1|m1@2 net264 i32|i0|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i1|i1|m1@2 net263 i32|i1|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i2|i1|m1@2 net262 i32|i2|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi32|i3|i1|m1@2 net261 i32|i3|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i0|i0|m1 i40|i0|net4 net229 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i0|i0|m1@2 i40|i0|net4 net229 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i0|i1|m1 q<3> i40|i0|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i0|i1|m1@2 q<3> i40|i0|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i1|i0|m1 i40|i1|net4 net227 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i1|i0|m1@2 i40|i1|net4 net227 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i1|i1|m1 q<2> i40|i1|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i1|i1|m1@2 q<2> i40|i1|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i2|i0|m1 i40|i2|net4 net225 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i2|i0|m1@2 i40|i2|net4 net225 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i2|i1|m1 q<1> i40|i2|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i2|i1|m1@2 q<1> i40|i2|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i3|i0|m1 i40|i3|net4 net355 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i3|i0|m1@2 i40|i3|net4 net355 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i3|i1|m1 q<0> i40|i3|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
mi40|i3|i1|m1@2 q<0> i40|i3|net4 vdd! pfet nfin=4 w=0.021u l=0.015u adeo=1.134e-15
+  aseo=5.67e-16 pdeo=2.34e-07 pseo=1.17e-07
cg662_5 i0|i57|i3|q 0  c=2.09084e-17
c662_4 i0|i57|i3|q i0|i59|i3|q  c=3.56053e-18
c662_3 i0|i57|i3|q i0|i57|i3|qb  c=3.06828e-17
c662_2 i0|i57|i3|q i0|i55|i3|q  c=4.07592e-18
c662_1 i0|i57|i3|q net263  c=1.27735e-17
cg661_5 i0|i57|i2|qb 0  c=2.98896e-17
c661_4 i0|i57|i2|qb i0|i57|i2|q  c=3.07268e-17
c661_3 i0|i57|i2|qb i0|i59|i2|qb  c=3.55906e-18
c661_2 i0|i57|i2|qb i0|i55|i2|qb  c=5.20112e-18
c661_1 i0|i57|i2|qb net263  c=5.82667e-18
cg660_4 i0|i57|i2|q 0  c=2.09006e-17
c660_3 i0|i57|i2|q i0|i59|i2|q  c=3.56053e-18
c660_2 i0|i57|i2|q i0|i55|i2|q  c=4.07592e-18
c660_1 i0|i57|i2|q net263  c=1.27789e-17
cg659_5 i0|i57|i1|qb 0  c=3.00078e-17
c659_4 i0|i57|i1|qb i0|i57|i1|q  c=3.06805e-17
c659_3 i0|i57|i1|qb i0|i59|i1|qb  c=3.55906e-18
c659_2 i0|i57|i1|qb i0|i55|i1|qb  c=5.20066e-18
c659_1 i0|i57|i1|qb net263  c=5.87913e-18
cg658_4 i0|i57|i1|q 0  c=2.0948e-17
c658_3 i0|i57|i1|q i0|i59|i1|q  c=3.56053e-18
c658_2 i0|i57|i1|q i0|i55|i1|q  c=4.07592e-18
c658_1 i0|i57|i1|q net263  c=1.26892e-17
cg657_5 i0|i57|i0|qb 0  c=2.99272e-17
c657_4 i0|i57|i0|qb i0|i57|i0|q  c=3.06656e-17
c657_3 i0|i57|i0|qb i0|i59|i0|qb  c=3.55906e-18
c657_2 i0|i57|i0|qb i0|i55|i0|qb  c=5.19742e-18
c657_1 i0|i57|i0|qb net263  c=5.79711e-18
cg656_4 i0|i57|i0|q 0  c=2.11391e-17
c656_3 i0|i57|i0|q i0|i59|i0|q  c=3.56053e-18
c656_2 i0|i57|i0|q i0|i55|i0|q  c=4.06641e-18
c656_1 i0|i57|i0|q net263  c=1.27286e-17
cg655_5 i0|i59|i3|qb 0  c=2.97975e-17
c655_4 i0|i59|i3|qb i0|i59|i3|q  c=3.07639e-17
c655_3 i0|i59|i3|qb i0|i57|i3|qb  c=3.55906e-18
c655_2 i0|i59|i3|qb i0|i61|i3|qb  c=5.20579e-18
c655_1 i0|i59|i3|qb net262  c=6.16568e-18
cg654_3 i0|i59|i3|q 0  c=2.14022e-17
c654_2 i0|i59|i3|q i0|i61|i3|q  c=4.07592e-18
c654_1 i0|i59|i3|q net262  c=1.20933e-17
cg653_4 i0|i59|i2|qb 0  c=2.9855e-17
c653_3 i0|i59|i2|qb i0|i59|i2|q  c=3.08127e-17
c653_2 i0|i59|i2|qb i0|i61|i2|qb  c=5.20112e-18
c653_1 i0|i59|i2|qb net262  c=6.02086e-18
cg652_3 i0|i59|i2|q 0  c=2.14014e-17
c652_2 i0|i59|i2|q i0|i61|i2|q  c=4.07592e-18
c652_1 i0|i59|i2|q net262  c=1.20954e-17
cg651_4 i0|i59|i1|qb 0  c=2.97956e-17
c651_3 i0|i59|i1|qb i0|i59|i1|q  c=3.07645e-17
c651_2 i0|i59|i1|qb i0|i61|i1|qb  c=5.20066e-18
c651_1 i0|i59|i1|qb net262  c=6.11153e-18
cg650_3 i0|i59|i1|q 0  c=2.14086e-17
c650_2 i0|i59|i1|q i0|i61|i1|q  c=4.07592e-18
c650_1 i0|i59|i1|q net262  c=1.20619e-17
cg649_4 i0|i59|i0|qb 0  c=2.9901e-17
c649_3 i0|i59|i0|qb i0|i59|i0|q  c=3.07502e-17
c649_2 i0|i59|i0|qb i0|i61|i0|qb  c=5.19742e-18
c649_1 i0|i59|i0|qb net262  c=6.06694e-18
cg648_3 i0|i59|i0|q 0  c=2.17107e-17
c648_2 i0|i59|i0|q i0|i61|i0|q  c=4.06641e-18
c648_1 i0|i59|i0|q net262  c=1.20572e-17
cg647_3 i0|i57|i3|qb 0  c=2.9935e-17
c647_2 i0|i57|i3|qb i0|i55|i3|qb  c=5.20579e-18
c647_1 i0|i57|i3|qb net263  c=5.89724e-18
cg614_5 i0|i49|i3|q 0  c=2.09061e-17
c614_4 i0|i49|i3|q i0|i51|i3|q  c=3.56053e-18
c614_3 i0|i49|i3|q i0|i49|i3|qb  c=3.06828e-17
c614_2 i0|i49|i3|q i0|i47|i3|q  c=4.07592e-18
c614_1 i0|i49|i3|q net271  c=1.27735e-17
cg613_5 i0|i49|i2|qb 0  c=2.9889e-17
c613_4 i0|i49|i2|qb i0|i49|i2|q  c=3.07268e-17
c613_3 i0|i49|i2|qb i0|i51|i2|qb  c=3.55906e-18
c613_2 i0|i49|i2|qb i0|i47|i2|qb  c=5.20112e-18
c613_1 i0|i49|i2|qb net271  c=5.82667e-18
cg612_4 i0|i49|i2|q 0  c=2.08984e-17
c612_3 i0|i49|i2|q i0|i51|i2|q  c=3.56053e-18
c612_2 i0|i49|i2|q i0|i47|i2|q  c=4.07592e-18
c612_1 i0|i49|i2|q net271  c=1.27789e-17
cg611_5 i0|i49|i1|qb 0  c=3.00072e-17
c611_4 i0|i49|i1|qb i0|i49|i1|q  c=3.06805e-17
c611_3 i0|i49|i1|qb i0|i51|i1|qb  c=3.55906e-18
c611_2 i0|i49|i1|qb i0|i47|i1|qb  c=5.20066e-18
c611_1 i0|i49|i1|qb net271  c=5.87913e-18
cg610_4 i0|i49|i1|q 0  c=2.09458e-17
c610_3 i0|i49|i1|q i0|i51|i1|q  c=3.56053e-18
c610_2 i0|i49|i1|q i0|i47|i1|q  c=4.07592e-18
c610_1 i0|i49|i1|q net271  c=1.26892e-17
cg609_5 i0|i49|i0|qb 0  c=2.99266e-17
c609_4 i0|i49|i0|qb i0|i49|i0|q  c=3.06656e-17
c609_3 i0|i49|i0|qb i0|i51|i0|qb  c=3.55906e-18
c609_2 i0|i49|i0|qb i0|i47|i0|qb  c=5.19742e-18
c609_1 i0|i49|i0|qb net271  c=5.79711e-18
cg608_4 i0|i49|i0|q 0  c=2.11368e-17
c608_3 i0|i49|i0|q i0|i51|i0|q  c=3.56053e-18
c608_2 i0|i49|i0|q i0|i47|i0|q  c=4.06641e-18
c608_1 i0|i49|i0|q net271  c=1.27286e-17
cg607_5 i0|i51|i3|qb 0  c=2.97775e-17
c607_4 i0|i51|i3|qb i0|i51|i3|q  c=3.07638e-17
c607_3 i0|i51|i3|qb i0|i49|i3|qb  c=3.55906e-18
c607_2 i0|i51|i3|qb i0|i53|i3|qb  c=5.20579e-18
c607_1 i0|i51|i3|qb net270  c=6.16568e-18
cg606_3 i0|i51|i3|q 0  c=2.13733e-17
c606_2 i0|i51|i3|q i0|i53|i3|q  c=4.07592e-18
c606_1 i0|i51|i3|q net270  c=1.20933e-17
cg605_4 i0|i51|i2|qb 0  c=2.9835e-17
c605_3 i0|i51|i2|qb i0|i51|i2|q  c=3.08125e-17
c605_2 i0|i51|i2|qb i0|i53|i2|qb  c=5.20112e-18
c605_1 i0|i51|i2|qb net270  c=6.02086e-18
cg604_3 i0|i51|i2|q 0  c=2.13726e-17
c604_2 i0|i51|i2|q i0|i53|i2|q  c=4.07592e-18
c604_1 i0|i51|i2|q net270  c=1.20954e-17
cg603_4 i0|i51|i1|qb 0  c=2.97761e-17
c603_3 i0|i51|i1|qb i0|i51|i1|q  c=3.07644e-17
c603_2 i0|i51|i1|qb i0|i53|i1|qb  c=5.20066e-18
c603_1 i0|i51|i1|qb net270  c=6.11153e-18
cg602_3 i0|i51|i1|q 0  c=2.13965e-17
c602_2 i0|i51|i1|q i0|i53|i1|q  c=4.07592e-18
c602_1 i0|i51|i1|q net270  c=1.20619e-17
cg601_4 i0|i51|i0|qb 0  c=2.98811e-17
c601_3 i0|i51|i0|qb i0|i51|i0|q  c=3.07499e-17
c601_2 i0|i51|i0|qb i0|i53|i0|qb  c=5.19742e-18
c601_1 i0|i51|i0|qb net270  c=6.06694e-18
cg600_3 i0|i51|i0|q 0  c=2.16817e-17
c600_2 i0|i51|i0|q i0|i53|i0|q  c=4.06641e-18
c600_1 i0|i51|i0|q net270  c=1.20572e-17
cg599_3 i0|i49|i3|qb 0  c=2.99344e-17
c599_2 i0|i49|i3|qb i0|i47|i3|qb  c=5.20579e-18
c599_1 i0|i49|i3|qb net271  c=5.89724e-18
cg566_5 i0|i41|i3|q 0  c=2.09027e-17
c566_4 i0|i41|i3|q i0|i43|i3|q  c=3.56053e-18
c566_3 i0|i41|i3|q i0|i41|i3|qb  c=3.06815e-17
c566_2 i0|i41|i3|q i0|i39|i3|q  c=4.07592e-18
c566_1 i0|i41|i3|q net275  c=1.27735e-17
cg565_5 i0|i41|i2|qb 0  c=2.9889e-17
c565_4 i0|i41|i2|qb i0|i41|i2|q  c=3.07255e-17
c565_3 i0|i41|i2|qb i0|i43|i2|qb  c=3.55906e-18
c565_2 i0|i41|i2|qb i0|i39|i2|qb  c=5.20112e-18
c565_1 i0|i41|i2|qb net275  c=5.82667e-18
cg564_4 i0|i41|i2|q 0  c=2.08949e-17
c564_3 i0|i41|i2|q i0|i43|i2|q  c=3.56053e-18
c564_2 i0|i41|i2|q i0|i39|i2|q  c=4.07592e-18
c564_1 i0|i41|i2|q net275  c=1.27789e-17
cg563_5 i0|i41|i1|qb 0  c=3.00071e-17
c563_4 i0|i41|i1|qb i0|i41|i1|q  c=3.06792e-17
c563_3 i0|i41|i1|qb i0|i43|i1|qb  c=3.55906e-18
c563_2 i0|i41|i1|qb i0|i39|i1|qb  c=5.20066e-18
c563_1 i0|i41|i1|qb net275  c=5.87913e-18
cg562_4 i0|i41|i1|q 0  c=2.09423e-17
c562_3 i0|i41|i1|q i0|i43|i1|q  c=3.56053e-18
c562_2 i0|i41|i1|q i0|i39|i1|q  c=4.07592e-18
c562_1 i0|i41|i1|q net275  c=1.26892e-17
cg561_5 i0|i41|i0|qb 0  c=2.99266e-17
c561_4 i0|i41|i0|qb i0|i41|i0|q  c=3.06643e-17
c561_3 i0|i41|i0|qb i0|i43|i0|qb  c=3.55906e-18
c561_2 i0|i41|i0|qb i0|i39|i0|qb  c=5.19742e-18
c561_1 i0|i41|i0|qb net275  c=5.79711e-18
cg560_4 i0|i41|i0|q 0  c=2.11333e-17
c560_3 i0|i41|i0|q i0|i43|i0|q  c=3.56053e-18
c560_2 i0|i41|i0|q i0|i39|i0|q  c=4.06641e-18
c560_1 i0|i41|i0|q net275  c=1.27286e-17
cg559_5 i0|i43|i3|qb 0  c=2.97637e-17
c559_4 i0|i43|i3|qb i0|i43|i3|q  c=3.07639e-17
c559_3 i0|i43|i3|qb i0|i41|i3|qb  c=3.55906e-18
c559_2 i0|i43|i3|qb i0|i45|i3|qb  c=5.20579e-18
c559_1 i0|i43|i3|qb net274  c=6.16624e-18
cg558_3 i0|i43|i3|q 0  c=2.13889e-17
c558_2 i0|i43|i3|q i0|i45|i3|q  c=4.07592e-18
c558_1 i0|i43|i3|q net274  c=1.20936e-17
cg557_4 i0|i43|i2|qb 0  c=2.98212e-17
c557_3 i0|i43|i2|qb i0|i43|i2|q  c=3.08127e-17
c557_2 i0|i43|i2|qb i0|i45|i2|qb  c=5.20112e-18
c557_1 i0|i43|i2|qb net274  c=6.02142e-18
cg556_3 i0|i43|i2|q 0  c=2.13882e-17
c556_2 i0|i43|i2|q i0|i45|i2|q  c=4.07592e-18
c556_1 i0|i43|i2|q net274  c=1.20957e-17
cg555_4 i0|i43|i1|qb 0  c=2.97618e-17
c555_3 i0|i43|i1|qb i0|i43|i1|q  c=3.07645e-17
c555_2 i0|i43|i1|qb i0|i45|i1|qb  c=5.20066e-18
c555_1 i0|i43|i1|qb net274  c=6.11209e-18
cg554_3 i0|i43|i1|q 0  c=2.14115e-17
c554_2 i0|i43|i1|q i0|i45|i1|q  c=4.07592e-18
c554_1 i0|i43|i1|q net274  c=1.20622e-17
cg553_4 i0|i43|i0|qb 0  c=2.98671e-17
c553_3 i0|i43|i0|qb i0|i43|i0|q  c=3.07502e-17
c553_2 i0|i43|i0|qb i0|i45|i0|qb  c=5.19742e-18
c553_1 i0|i43|i0|qb net274  c=6.0675e-18
cg552_3 i0|i43|i0|q 0  c=2.16828e-17
c552_2 i0|i43|i0|q i0|i45|i0|q  c=4.06641e-18
c552_1 i0|i43|i0|q net274  c=1.20575e-17
cg551_3 i0|i41|i3|qb 0  c=2.99344e-17
c551_2 i0|i41|i3|qb i0|i39|i3|qb  c=5.20579e-18
c551_1 i0|i41|i3|qb net275  c=5.89724e-18
cg518_5 i0|i33|i3|q 0  c=2.09145e-17
c518_4 i0|i33|i3|q i0|i35|i3|q  c=3.56053e-18
c518_3 i0|i33|i3|q i0|i33|i3|qb  c=3.06828e-17
c518_2 i0|i33|i3|q i0|i31|i3|q  c=4.07592e-18
c518_1 i0|i33|i3|q net279  c=1.27735e-17
cg517_5 i0|i33|i2|qb 0  c=2.99039e-17
c517_4 i0|i33|i2|qb i0|i33|i2|q  c=3.07268e-17
c517_3 i0|i33|i2|qb i0|i35|i2|qb  c=3.55906e-18
c517_2 i0|i33|i2|qb i0|i31|i2|qb  c=5.20112e-18
c517_1 i0|i33|i2|qb net279  c=5.82667e-18
cg516_4 i0|i33|i2|q 0  c=2.0918e-17
c516_3 i0|i33|i2|q i0|i35|i2|q  c=3.56053e-18
c516_2 i0|i33|i2|q i0|i31|i2|q  c=4.07592e-18
c516_1 i0|i33|i2|q net279  c=1.25763e-17
cg515_5 i0|i33|i1|qb 0  c=2.99346e-17
c515_4 i0|i33|i1|qb i0|i33|i1|q  c=3.06805e-17
c515_3 i0|i33|i1|qb i0|i35|i1|qb  c=3.55906e-18
c515_2 i0|i33|i1|qb i0|i31|i1|qb  c=5.18719e-18
c515_1 i0|i33|i1|qb net279  c=5.87913e-18
cg514_4 i0|i33|i1|q 0  c=2.09479e-17
c514_3 i0|i33|i1|q i0|i35|i1|q  c=3.56053e-18
c514_2 i0|i33|i1|q i0|i31|i1|q  c=4.07592e-18
c514_1 i0|i33|i1|q net279  c=1.26892e-17
cg513_5 i0|i33|i0|qb 0  c=2.99415e-17
c513_4 i0|i33|i0|qb i0|i33|i0|q  c=3.06656e-17
c513_3 i0|i33|i0|qb i0|i35|i0|qb  c=3.55906e-18
c513_2 i0|i33|i0|qb i0|i31|i0|qb  c=5.19742e-18
c513_1 i0|i33|i0|qb net279  c=5.79711e-18
cg512_4 i0|i33|i0|q 0  c=2.11564e-17
c512_3 i0|i33|i0|q i0|i35|i0|q  c=3.56053e-18
c512_2 i0|i33|i0|q i0|i31|i0|q  c=4.06641e-18
c512_1 i0|i33|i0|q net279  c=1.25271e-17
cg511_5 i0|i35|i3|qb 0  c=2.97777e-17
c511_4 i0|i35|i3|qb i0|i35|i3|q  c=3.07639e-17
c511_3 i0|i35|i3|qb i0|i33|i3|qb  c=3.55906e-18
c511_2 i0|i35|i3|qb i0|i37|i3|qb  c=5.20579e-18
c511_1 i0|i35|i3|qb net278  c=6.16568e-18
cg510_3 i0|i35|i3|q 0  c=2.13748e-17
c510_2 i0|i35|i3|q i0|i37|i3|q  c=4.07592e-18
c510_1 i0|i35|i3|q net278  c=1.20933e-17
cg509_4 i0|i35|i2|qb 0  c=2.98352e-17
c509_3 i0|i35|i2|qb i0|i35|i2|q  c=3.08127e-17
c509_2 i0|i35|i2|qb i0|i37|i2|qb  c=5.20112e-18
c509_1 i0|i35|i2|qb net278  c=6.02086e-18
cg508_3 i0|i35|i2|q 0  c=2.1374e-17
c508_2 i0|i35|i2|q i0|i37|i2|q  c=4.07592e-18
c508_1 i0|i35|i2|q net278  c=1.20954e-17
cg507_4 i0|i35|i1|qb 0  c=2.97758e-17
c507_3 i0|i35|i1|qb i0|i35|i1|q  c=3.07645e-17
c507_2 i0|i35|i1|qb i0|i37|i1|qb  c=5.20066e-18
c507_1 i0|i35|i1|qb net278  c=6.11153e-18
cg506_3 i0|i35|i1|q 0  c=2.13971e-17
c506_2 i0|i35|i1|q i0|i37|i1|q  c=4.07592e-18
c506_1 i0|i35|i1|q net278  c=1.20619e-17
cg505_4 i0|i35|i0|qb 0  c=2.98811e-17
c505_3 i0|i35|i0|qb i0|i35|i0|q  c=3.07502e-17
c505_2 i0|i35|i0|qb i0|i37|i0|qb  c=5.19742e-18
c505_1 i0|i35|i0|qb net278  c=6.06694e-18
cg504_3 i0|i35|i0|q 0  c=2.16834e-17
c504_2 i0|i35|i0|q i0|i37|i0|q  c=4.06641e-18
c504_1 i0|i35|i0|q net278  c=1.20572e-17
cg503_3 i0|i33|i3|qb 0  c=2.99295e-17
c503_2 i0|i33|i3|qb i0|i31|i3|qb  c=5.20579e-18
c503_1 i0|i33|i3|qb net279  c=5.89724e-18
cg470_5 i0|i56|i3|q 0  c=2.06501e-17
c470_4 i0|i56|i3|q i0|i58|i3|q  c=3.56162e-18
c470_3 i0|i56|i3|q i0|i56|i3|qb  c=3.0708e-17
c470_2 i0|i56|i3|q i0|i54|i3|q  c=4.07691e-18
c470_1 i0|i56|i3|q net263  c=1.29968e-17
cg469_5 i0|i56|i2|qb 0  c=3.00159e-17
c469_4 i0|i56|i2|qb i0|i56|i2|q  c=3.06805e-17
c469_3 i0|i56|i2|qb i0|i58|i2|qb  c=3.55906e-18
c469_2 i0|i56|i2|qb i0|i54|i2|qb  c=5.20066e-18
c469_1 i0|i56|i2|qb net263  c=5.88004e-18
cg468_4 i0|i56|i2|q 0  c=2.09307e-17
c468_3 i0|i56|i2|q i0|i58|i2|q  c=3.56053e-18
c468_2 i0|i56|i2|q i0|i54|i2|q  c=4.07592e-18
c468_1 i0|i56|i2|q net263  c=1.27096e-17
cg467_5 i0|i56|i1|qb 0  c=2.99028e-17
c467_4 i0|i56|i1|qb i0|i56|i1|q  c=3.07268e-17
c467_3 i0|i56|i1|qb i0|i58|i1|qb  c=3.55906e-18
c467_2 i0|i56|i1|qb i0|i54|i1|qb  c=5.19742e-18
c467_1 i0|i56|i1|qb net263  c=5.79874e-18
cg466_4 i0|i56|i1|q 0  c=2.08972e-17
c466_3 i0|i56|i1|q i0|i58|i1|q  c=3.56053e-18
c466_2 i0|i56|i1|q i0|i54|i1|q  c=4.07592e-18
c466_1 i0|i56|i1|q net263  c=1.27792e-17
cg465_5 i0|i56|i0|qb 0  c=3.00619e-17
c465_4 i0|i56|i0|qb i0|i56|i0|q  c=3.06823e-17
c465_3 i0|i56|i0|qb i0|i58|i0|qb  c=3.55906e-18
c465_2 i0|i56|i0|qb i0|i54|i0|qb  c=5.19561e-18
c465_1 i0|i56|i0|qb net263  c=5.86113e-18
cg464_4 i0|i56|i0|q 0  c=2.1057e-17
c464_3 i0|i56|i0|q i0|i58|i0|q  c=3.56053e-18
c464_2 i0|i56|i0|q i0|i54|i0|q  c=4.06766e-18
c464_1 i0|i56|i0|q net263  c=1.26447e-17
cg463_5 i0|i58|i3|qb 0  c=2.96557e-17
c463_4 i0|i58|i3|qb i0|i58|i3|q  c=3.07503e-17
c463_3 i0|i58|i3|qb i0|i56|i3|qb  c=3.55906e-18
c463_2 i0|i58|i3|qb i0|i60|i3|qb  c=5.20112e-18
c463_1 i0|i58|i3|qb net262  c=6.08559e-18
cg462_3 i0|i58|i3|q 0  c=2.09641e-17
c462_2 i0|i58|i3|q i0|i60|i3|q  c=4.07691e-18
c462_1 i0|i58|i3|q net262  c=1.23905e-17
cg461_4 i0|i58|i2|qb 0  c=2.98807e-17
c461_3 i0|i58|i2|qb i0|i58|i2|q  c=3.07667e-17
c461_2 i0|i58|i2|qb i0|i60|i2|qb  c=5.20066e-18
c461_1 i0|i58|i2|qb net262  c=6.10567e-18
cg460_3 i0|i58|i2|q 0  c=2.14087e-17
c460_2 i0|i58|i2|q i0|i60|i2|q  c=4.07592e-18
c460_1 i0|i58|i2|q net262  c=1.20747e-17
cg459_4 i0|i58|i1|qb 0  c=2.98566e-17
c459_3 i0|i58|i1|qb i0|i58|i1|q  c=3.08127e-17
c459_2 i0|i58|i1|qb i0|i60|i1|qb  c=5.19742e-18
c459_1 i0|i58|i1|qb net262  c=6.01587e-18
cg458_3 i0|i58|i1|q 0  c=2.1407e-17
c458_2 i0|i58|i1|q i0|i60|i1|q  c=4.07592e-18
c458_1 i0|i58|i1|q net262  c=1.20928e-17
cg457_4 i0|i58|i0|qb 0  c=2.99145e-17
c457_3 i0|i58|i0|qb i0|i58|i0|q  c=3.07592e-17
c457_2 i0|i58|i0|qb i0|i60|i0|qb  c=5.19561e-18
c457_1 i0|i58|i0|qb net262  c=6.14999e-18
cg456_3 i0|i58|i0|q 0  c=2.1475e-17
c456_2 i0|i58|i0|q i0|i60|i0|q  c=4.06766e-18
c456_1 i0|i58|i0|q net262  c=1.20485e-17
cg455_3 i0|i56|i3|qb 0  c=2.97014e-17
c455_2 i0|i56|i3|qb i0|i54|i3|qb  c=5.20112e-18
c455_1 i0|i56|i3|qb net263  c=5.99239e-18
cg422_5 i0|i48|i3|q 0  c=2.06222e-17
c422_4 i0|i48|i3|q i0|i50|i3|q  c=3.56162e-18
c422_3 i0|i48|i3|q i0|i48|i3|qb  c=3.0708e-17
c422_2 i0|i48|i3|q i0|i46|i3|q  c=4.07691e-18
c422_1 i0|i48|i3|q net271  c=1.29968e-17
cg421_5 i0|i48|i2|qb 0  c=3.00153e-17
c421_4 i0|i48|i2|qb i0|i48|i2|q  c=3.06805e-17
c421_3 i0|i48|i2|qb i0|i50|i2|qb  c=3.55906e-18
c421_2 i0|i48|i2|qb i0|i46|i2|qb  c=5.20066e-18
c421_1 i0|i48|i2|qb net271  c=5.88004e-18
cg420_4 i0|i48|i2|q 0  c=2.09284e-17
c420_3 i0|i48|i2|q i0|i50|i2|q  c=3.56053e-18
c420_2 i0|i48|i2|q i0|i46|i2|q  c=4.07592e-18
c420_1 i0|i48|i2|q net271  c=1.27096e-17
cg419_5 i0|i48|i1|qb 0  c=2.99021e-17
c419_4 i0|i48|i1|qb i0|i48|i1|q  c=3.07268e-17
c419_3 i0|i48|i1|qb i0|i50|i1|qb  c=3.55906e-18
c419_2 i0|i48|i1|qb i0|i46|i1|qb  c=5.19742e-18
c419_1 i0|i48|i1|qb net271  c=5.79874e-18
cg418_4 i0|i48|i1|q 0  c=2.08949e-17
c418_3 i0|i48|i1|q i0|i50|i1|q  c=3.56053e-18
c418_2 i0|i48|i1|q i0|i46|i1|q  c=4.07592e-18
c418_1 i0|i48|i1|q net271  c=1.27792e-17
cg417_5 i0|i48|i0|qb 0  c=3.00613e-17
c417_4 i0|i48|i0|qb i0|i48|i0|q  c=3.06823e-17
c417_3 i0|i48|i0|qb i0|i50|i0|qb  c=3.55906e-18
c417_2 i0|i48|i0|qb i0|i46|i0|qb  c=5.19561e-18
c417_1 i0|i48|i0|qb net271  c=5.86113e-18
cg416_4 i0|i48|i0|q 0  c=2.10547e-17
c416_3 i0|i48|i0|q i0|i50|i0|q  c=3.56053e-18
c416_2 i0|i48|i0|q i0|i46|i0|q  c=4.06766e-18
c416_1 i0|i48|i0|q net271  c=1.26447e-17
cg415_5 i0|i50|i3|qb 0  c=2.96383e-17
c415_4 i0|i50|i3|qb i0|i50|i3|q  c=3.07501e-17
c415_3 i0|i50|i3|qb i0|i48|i3|qb  c=3.55906e-18
c415_2 i0|i50|i3|qb i0|i52|i3|qb  c=5.20112e-18
c415_1 i0|i50|i3|qb net270  c=6.08559e-18
cg414_3 i0|i50|i3|q 0  c=2.09366e-17
c414_2 i0|i50|i3|q i0|i52|i3|q  c=4.07691e-18
c414_1 i0|i50|i3|q net270  c=1.23905e-17
cg413_4 i0|i50|i2|qb 0  c=2.98608e-17
c413_3 i0|i50|i2|qb i0|i50|i2|q  c=3.07665e-17
c413_2 i0|i50|i2|qb i0|i52|i2|qb  c=5.20066e-18
c413_1 i0|i50|i2|qb net270  c=6.10567e-18
cg412_3 i0|i50|i2|q 0  c=2.13798e-17
c412_2 i0|i50|i2|q i0|i52|i2|q  c=4.07592e-18
c412_1 i0|i50|i2|q net270  c=1.20747e-17
cg411_4 i0|i50|i1|qb 0  c=2.98367e-17
c411_3 i0|i50|i1|qb i0|i50|i1|q  c=3.08125e-17
c411_2 i0|i50|i1|qb i0|i52|i1|qb  c=5.19742e-18
c411_1 i0|i50|i1|qb net270  c=6.01587e-18
cg410_3 i0|i50|i1|q 0  c=2.13781e-17
c410_2 i0|i50|i1|q i0|i52|i1|q  c=4.07592e-18
c410_1 i0|i50|i1|q net270  c=1.20928e-17
cg409_4 i0|i50|i0|qb 0  c=2.98944e-17
c409_3 i0|i50|i0|qb i0|i50|i0|q  c=3.0759e-17
c409_2 i0|i50|i0|qb i0|i52|i0|qb  c=5.19561e-18
c409_1 i0|i50|i0|qb net270  c=6.14999e-18
cg408_3 i0|i50|i0|q 0  c=2.14902e-17
c408_2 i0|i50|i0|q i0|i52|i0|q  c=4.06766e-18
c408_1 i0|i50|i0|q net270  c=1.20485e-17
cg407_3 i0|i48|i3|qb 0  c=2.97014e-17
c407_2 i0|i48|i3|qb i0|i46|i3|qb  c=5.20112e-18
c407_1 i0|i48|i3|qb net271  c=5.99239e-18
cg374_5 i0|i40|i3|q 0  c=2.06187e-17
c374_4 i0|i40|i3|q i0|i42|i3|q  c=3.56162e-18
c374_3 i0|i40|i3|q i0|i40|i3|qb  c=3.07067e-17
c374_2 i0|i40|i3|q i0|i38|i3|q  c=4.07691e-18
c374_1 i0|i40|i3|q net275  c=1.29959e-17
cg373_5 i0|i40|i2|qb 0  c=3.00153e-17
c373_4 i0|i40|i2|qb i0|i40|i2|q  c=3.06792e-17
c373_3 i0|i40|i2|qb i0|i42|i2|qb  c=3.55906e-18
c373_2 i0|i40|i2|qb i0|i38|i2|qb  c=5.20066e-18
c373_1 i0|i40|i2|qb net275  c=5.88004e-18
cg372_4 i0|i40|i2|q 0  c=2.0925e-17
c372_3 i0|i40|i2|q i0|i42|i2|q  c=3.56053e-18
c372_2 i0|i40|i2|q i0|i38|i2|q  c=4.07592e-18
c372_1 i0|i40|i2|q net275  c=1.27096e-17
cg371_5 i0|i40|i1|qb 0  c=2.99021e-17
c371_4 i0|i40|i1|qb i0|i40|i1|q  c=3.07255e-17
c371_3 i0|i40|i1|qb i0|i42|i1|qb  c=3.55906e-18
c371_2 i0|i40|i1|qb i0|i38|i1|qb  c=5.19742e-18
c371_1 i0|i40|i1|qb net275  c=5.79874e-18
cg370_4 i0|i40|i1|q 0  c=2.08915e-17
c370_3 i0|i40|i1|q i0|i42|i1|q  c=3.56053e-18
c370_2 i0|i40|i1|q i0|i38|i1|q  c=4.07592e-18
c370_1 i0|i40|i1|q net275  c=1.27792e-17
cg369_5 i0|i40|i0|qb 0  c=3.00613e-17
c369_4 i0|i40|i0|qb i0|i40|i0|q  c=3.0681e-17
c369_3 i0|i40|i0|qb i0|i42|i0|qb  c=3.55906e-18
c369_2 i0|i40|i0|qb i0|i38|i0|qb  c=5.19561e-18
c369_1 i0|i40|i0|qb net275  c=5.86113e-18
cg368_4 i0|i40|i0|q 0  c=2.10513e-17
c368_3 i0|i40|i0|q i0|i42|i0|q  c=3.56053e-18
c368_2 i0|i40|i0|q i0|i38|i0|q  c=4.06766e-18
c368_1 i0|i40|i0|q net275  c=1.26447e-17
cg367_5 i0|i42|i3|qb 0  c=2.96385e-17
c367_4 i0|i42|i3|qb i0|i42|i3|q  c=3.07503e-17
c367_3 i0|i42|i3|qb i0|i40|i3|qb  c=3.55906e-18
c367_2 i0|i42|i3|qb i0|i44|i3|qb  c=5.20112e-18
c367_1 i0|i42|i3|qb net274  c=6.08381e-18
cg366_3 i0|i42|i3|q 0  c=2.09515e-17
c366_2 i0|i42|i3|q i0|i44|i3|q  c=4.07691e-18
c366_1 i0|i42|i3|q net274  c=1.23908e-17
cg365_4 i0|i42|i2|qb 0  c=2.98469e-17
c365_3 i0|i42|i2|qb i0|i42|i2|q  c=3.07667e-17
c365_2 i0|i42|i2|qb i0|i44|i2|qb  c=5.20066e-18
c365_1 i0|i42|i2|qb net274  c=6.10654e-18
cg364_3 i0|i42|i2|q 0  c=2.13954e-17
c364_2 i0|i42|i2|q i0|i44|i2|q  c=4.07592e-18
c364_1 i0|i42|i2|q net274  c=1.2075e-17
cg363_4 i0|i42|i1|qb 0  c=2.98229e-17
c363_3 i0|i42|i1|qb i0|i42|i1|q  c=3.08127e-17
c363_2 i0|i42|i1|qb i0|i44|i1|qb  c=5.19742e-18
c363_1 i0|i42|i1|qb net274  c=6.01674e-18
cg362_3 i0|i42|i1|q 0  c=2.13938e-17
c362_2 i0|i42|i1|q i0|i44|i1|q  c=4.07592e-18
c362_1 i0|i42|i1|q net274  c=1.20931e-17
cg361_4 i0|i42|i0|qb 0  c=2.98807e-17
c361_3 i0|i42|i0|qb i0|i42|i0|q  c=3.07592e-17
c361_2 i0|i42|i0|qb i0|i44|i0|qb  c=5.19561e-18
c361_1 i0|i42|i0|qb net274  c=6.15056e-18
cg360_3 i0|i42|i0|q 0  c=2.15054e-17
c360_2 i0|i42|i0|q i0|i44|i0|q  c=4.06766e-18
c360_1 i0|i42|i0|q net274  c=1.20488e-17
cg359_3 i0|i40|i3|qb 0  c=2.97047e-17
c359_2 i0|i40|i3|qb i0|i38|i3|qb  c=5.20112e-18
c359_1 i0|i40|i3|qb net275  c=5.99196e-18
cg326_5 i0|i32|i3|q 0  c=2.06421e-17
c326_4 i0|i32|i3|q i0|i34|i3|q  c=3.56162e-18
c326_3 i0|i32|i3|q i0|i32|i3|qb  c=3.0708e-17
c326_2 i0|i32|i3|q i0|i30|i3|q  c=4.07691e-18
c326_1 i0|i32|i3|q net279  c=1.28617e-17
cg325_5 i0|i32|i2|qb 0  c=2.9954e-17
c325_4 i0|i32|i2|qb i0|i32|i2|q  c=3.06805e-17
c325_3 i0|i32|i2|qb i0|i34|i2|qb  c=3.55906e-18
c325_2 i0|i32|i2|qb i0|i30|i2|qb  c=5.18719e-18
c325_1 i0|i32|i2|qb net279  c=5.88004e-18
cg324_4 i0|i32|i2|q 0  c=2.09418e-17
c324_3 i0|i32|i2|q i0|i34|i2|q  c=3.56053e-18
c324_2 i0|i32|i2|q i0|i30|i2|q  c=4.07592e-18
c324_1 i0|i32|i2|q net279  c=1.27096e-17
cg323_5 i0|i32|i1|qb 0  c=2.99059e-17
c323_4 i0|i32|i1|qb i0|i32|i1|q  c=3.07268e-17
c323_3 i0|i32|i1|qb i0|i34|i1|qb  c=3.55906e-18
c323_2 i0|i32|i1|qb i0|i30|i1|qb  c=5.19742e-18
c323_1 i0|i32|i1|qb net279  c=5.79874e-18
cg322_4 i0|i32|i1|q 0  c=2.09033e-17
c322_3 i0|i32|i1|q i0|i34|i1|q  c=3.56053e-18
c322_2 i0|i32|i1|q i0|i30|i1|q  c=4.07592e-18
c322_1 i0|i32|i1|q net279  c=1.27792e-17
cg321_5 i0|i32|i0|qb 0  c=3.00226e-17
c321_4 i0|i32|i0|qb i0|i32|i0|q  c=3.06823e-17
c321_3 i0|i32|i0|qb i0|i34|i0|qb  c=3.55906e-18
c321_2 i0|i32|i0|qb i0|i30|i0|qb  c=5.19561e-18
c321_1 i0|i32|i0|qb net279  c=5.86113e-18
cg320_4 i0|i32|i0|q 0  c=2.10655e-17
c320_3 i0|i32|i0|q i0|i34|i0|q  c=3.56053e-18
c320_2 i0|i32|i0|q i0|i30|i0|q  c=4.06766e-18
c320_1 i0|i32|i0|q net279  c=1.25259e-17
cg319_5 i0|i34|i3|qb 0  c=2.9637e-17
c319_4 i0|i34|i3|qb i0|i34|i3|q  c=3.07503e-17
c319_3 i0|i34|i3|qb i0|i32|i3|qb  c=3.55906e-18
c319_2 i0|i34|i3|qb i0|i36|i3|qb  c=5.20112e-18
c319_1 i0|i34|i3|qb net278  c=6.08301e-18
cg318_3 i0|i34|i3|q 0  c=2.09368e-17
c318_2 i0|i34|i3|q i0|i36|i3|q  c=4.07691e-18
c318_1 i0|i34|i3|q net278  c=1.23905e-17
cg317_4 i0|i34|i2|qb 0  c=2.98609e-17
c317_3 i0|i34|i2|qb i0|i34|i2|q  c=3.07667e-17
c317_2 i0|i34|i2|qb i0|i36|i2|qb  c=5.20066e-18
c317_1 i0|i34|i2|qb net278  c=6.10567e-18
cg316_3 i0|i34|i2|q 0  c=2.13814e-17
c316_2 i0|i34|i2|q i0|i36|i2|q  c=4.07592e-18
c316_1 i0|i34|i2|q net278  c=1.20747e-17
cg315_4 i0|i34|i1|qb 0  c=2.98369e-17
c315_3 i0|i34|i1|qb i0|i34|i1|q  c=3.08127e-17
c315_2 i0|i34|i1|qb i0|i36|i1|qb  c=5.19742e-18
c315_1 i0|i34|i1|qb net278  c=6.01587e-18
cg314_3 i0|i34|i1|q 0  c=2.13796e-17
c314_2 i0|i34|i1|q i0|i36|i1|q  c=4.07592e-18
c314_1 i0|i34|i1|q net278  c=1.20928e-17
cg313_4 i0|i34|i0|qb 0  c=2.98947e-17
c313_3 i0|i34|i0|qb i0|i34|i0|q  c=3.07592e-17
c313_2 i0|i34|i0|qb i0|i36|i0|qb  c=5.19561e-18
c313_1 i0|i34|i0|qb net278  c=6.14999e-18
cg312_3 i0|i34|i0|q 0  c=2.14911e-17
c312_2 i0|i34|i0|q i0|i36|i0|q  c=4.06766e-18
c312_1 i0|i34|i0|q net278  c=1.20485e-17
cg311_3 i0|i32|i3|qb 0  c=2.97191e-17
c311_2 i0|i32|i3|qb i0|i30|i3|qb  c=5.20112e-18
c311_1 i0|i32|i3|qb net279  c=5.99196e-18
cg310_4 i0|i45|i0|qb 0  c=2.99266e-17
c310_3 i0|i45|i0|qb i0|i45|i0|q  c=3.06656e-17
c310_2 i0|i45|i0|qb i0|i47|i0|qb  c=3.55906e-18
c310_1 i0|i45|i0|qb net273  c=5.79711e-18
cg309_3 i0|i45|i0|q 0  c=2.11368e-17
c309_2 i0|i45|i0|q i0|i47|i0|q  c=3.56053e-18
c309_1 i0|i45|i0|q net273  c=1.27286e-17
cg308_4 i0|i39|i3|qb 0  c=2.97777e-17
c308_3 i0|i39|i3|qb i0|i39|i3|q  c=3.07639e-17
c308_2 i0|i39|i3|qb i0|i37|i3|qb  c=3.55906e-18
c308_1 i0|i39|i3|qb net276  c=6.16568e-18
cg307_3 i0|i39|i3|q 0  c=2.13748e-17
c307_2 i0|i39|i3|q i0|i37|i3|q  c=3.56053e-18
c307_1 i0|i39|i3|q net276  c=1.20933e-17
cg306_4 i0|i39|i2|qb 0  c=2.98352e-17
c306_3 i0|i39|i2|qb i0|i39|i2|q  c=3.08127e-17
c306_2 i0|i39|i2|qb i0|i37|i2|qb  c=3.55906e-18
c306_1 i0|i39|i2|qb net276  c=6.02086e-18
cg305_3 i0|i39|i2|q 0  c=2.1374e-17
c305_2 i0|i39|i2|q i0|i37|i2|q  c=3.56053e-18
c305_1 i0|i39|i2|q net276  c=1.20954e-17
cg304_4 i0|i39|i1|qb 0  c=2.97758e-17
c304_3 i0|i39|i1|qb i0|i39|i1|q  c=3.07645e-17
c304_2 i0|i39|i1|qb i0|i37|i1|qb  c=3.55906e-18
c304_1 i0|i39|i1|qb net276  c=6.11153e-18
cg303_3 i0|i39|i1|q 0  c=2.13971e-17
c303_2 i0|i39|i1|q i0|i37|i1|q  c=3.56053e-18
c303_1 i0|i39|i1|q net276  c=1.20619e-17
cg302_4 i0|i39|i0|qb 0  c=2.98811e-17
c302_3 i0|i39|i0|qb i0|i39|i0|q  c=3.07502e-17
c302_2 i0|i39|i0|qb i0|i37|i0|qb  c=3.55906e-18
c302_1 i0|i39|i0|qb net276  c=6.06693e-18
cg301_3 i0|i39|i0|q 0  c=2.16834e-17
c301_2 i0|i39|i0|q i0|i37|i0|q  c=3.56053e-18
c301_1 i0|i39|i0|q net276  c=1.20572e-17
cg300_3 i0|i37|i3|qb 0  c=2.99344e-17
c300_2 i0|i37|i3|qb i0|i37|i3|q  c=3.06828e-17
c300_1 i0|i37|i3|qb net277  c=5.89724e-18
cg299_2 i0|i37|i3|q 0  c=2.09061e-17
c299_1 i0|i37|i3|q net277  c=1.27735e-17
cg298_3 i0|i37|i2|qb 0  c=2.9889e-17
c298_2 i0|i37|i2|qb i0|i37|i2|q  c=3.07268e-17
c298_1 i0|i37|i2|qb net277  c=5.82667e-18
cg297_2 i0|i37|i2|q 0  c=2.08984e-17
c297_1 i0|i37|i2|q net277  c=1.27789e-17
cg296_3 i0|i37|i1|qb 0  c=3.00072e-17
c296_2 i0|i37|i1|qb i0|i37|i1|q  c=3.06805e-17
c296_1 i0|i37|i1|qb net277  c=5.87913e-18
cg295_2 i0|i37|i1|q 0  c=2.09458e-17
c295_1 i0|i37|i1|q net277  c=1.26892e-17
cg294_3 i0|i37|i0|qb 0  c=2.99266e-17
c294_2 i0|i37|i0|qb i0|i37|i0|q  c=3.06656e-17
c294_1 i0|i37|i0|qb net277  c=5.79711e-18
cg293_2 i0|i37|i0|q 0  c=2.11368e-17
c293_1 i0|i37|i0|q net277  c=1.27286e-17
cg292_4 i0|i54|i3|qb 0  c=2.96405e-17
c292_3 i0|i54|i3|qb i0|i54|i3|q  c=3.07312e-17
c292_2 i0|i54|i3|qb i0|i52|i3|qb  c=3.55906e-18
c292_1 i0|i54|i3|qb net264  c=6.08559e-18
cg291_3 i0|i54|i3|q 0  c=2.09257e-17
c291_2 i0|i54|i3|q i0|i52|i3|q  c=3.56162e-18
c291_1 i0|i54|i3|q net264  c=1.23905e-17
cg290_4 i0|i54|i2|qb 0  c=2.98735e-17
c290_3 i0|i54|i2|qb i0|i54|i2|q  c=3.07512e-17
c290_2 i0|i54|i2|qb i0|i52|i2|qb  c=3.55906e-18
c290_1 i0|i54|i2|qb net264  c=6.10567e-18
cg289_3 i0|i54|i2|q 0  c=2.13935e-17
c289_2 i0|i54|i2|q i0|i52|i2|q  c=3.56053e-18
c289_1 i0|i54|i2|q net264  c=1.20747e-17
cg288_4 i0|i54|i1|qb 0  c=2.98494e-17
c288_3 i0|i54|i1|qb i0|i54|i1|q  c=3.07931e-17
c288_2 i0|i54|i1|qb i0|i52|i1|qb  c=3.55906e-18
c288_1 i0|i54|i1|qb net264  c=6.01587e-18
cg287_3 i0|i54|i1|q 0  c=2.13799e-17
c287_2 i0|i54|i1|q i0|i52|i1|q  c=3.56053e-18
c287_1 i0|i54|i1|q net264  c=1.20928e-17
cg286_4 i0|i54|i0|qb 0  c=2.99072e-17
c286_3 i0|i54|i0|qb i0|i54|i0|q  c=3.07437e-17
c286_2 i0|i54|i0|qb i0|i52|i0|qb  c=3.55906e-18
c286_1 i0|i54|i0|qb net264  c=6.14999e-18
cg285_3 i0|i54|i0|q 0  c=2.15081e-17
c285_2 i0|i54|i0|q i0|i52|i0|q  c=3.56053e-18
c285_1 i0|i54|i0|q net264  c=1.20485e-17
cg284_3 i0|i52|i3|qb 0  c=2.97021e-17
c284_2 i0|i52|i3|qb i0|i52|i3|q  c=3.0708e-17
c284_1 i0|i52|i3|qb net269  c=5.99239e-18
cg283_2 i0|i52|i3|q 0  c=2.06318e-17
c283_1 i0|i52|i3|q net269  c=1.29968e-17
cg282_3 i0|i52|i2|qb 0  c=3.00159e-17
c282_2 i0|i52|i2|qb i0|i52|i2|q  c=3.06805e-17
c282_1 i0|i52|i2|qb net269  c=5.88004e-18
cg281_2 i0|i52|i2|q 0  c=2.09271e-17
c281_1 i0|i52|i2|q net269  c=1.27058e-17
cg280_3 i0|i52|i1|qb 0  c=2.99028e-17
c280_2 i0|i52|i1|qb i0|i52|i1|q  c=3.07268e-17
c280_1 i0|i52|i1|qb net269  c=5.79874e-18
cg279_2 i0|i52|i1|q 0  c=2.08936e-17
c279_1 i0|i52|i1|q net269  c=1.27792e-17
cg278_3 i0|i52|i0|qb 0  c=3.00619e-17
c278_2 i0|i52|i0|qb i0|i52|i0|q  c=3.06823e-17
c278_1 i0|i52|i0|qb net269  c=5.86113e-18
cg277_2 i0|i52|i0|q 0  c=2.10534e-17
c277_1 i0|i52|i0|q net269  c=1.26421e-17
cg276_4 i0|i46|i3|qb 0  c=2.9639e-17
c276_3 i0|i46|i3|qb i0|i46|i3|q  c=3.07503e-17
c276_2 i0|i46|i3|qb i0|i44|i3|qb  c=3.55906e-18
c276_1 i0|i46|i3|qb net272  c=6.08559e-18
cg275_3 i0|i46|i3|q 0  c=2.09515e-17
c275_2 i0|i46|i3|q i0|i44|i3|q  c=3.56162e-18
c275_1 i0|i46|i3|q net272  c=1.23905e-17
cg274_4 i0|i46|i2|qb 0  c=2.98469e-17
c274_3 i0|i46|i2|qb i0|i46|i2|q  c=3.07667e-17
c274_2 i0|i46|i2|qb i0|i44|i2|qb  c=3.55906e-18
c274_1 i0|i46|i2|qb net272  c=6.10567e-18
cg273_3 i0|i46|i2|q 0  c=2.1395e-17
c273_2 i0|i46|i2|q i0|i44|i2|q  c=3.56053e-18
c273_1 i0|i46|i2|q net272  c=1.20747e-17
cg272_4 i0|i46|i1|qb 0  c=2.98229e-17
c272_3 i0|i46|i1|qb i0|i46|i1|q  c=3.08127e-17
c272_2 i0|i46|i1|qb i0|i44|i1|qb  c=3.55906e-18
c272_1 i0|i46|i1|qb net272  c=6.01587e-18
cg271_3 i0|i46|i1|q 0  c=2.13935e-17
c271_2 i0|i46|i1|q i0|i44|i1|q  c=3.56053e-18
c271_1 i0|i46|i1|q net272  c=1.20928e-17
cg270_4 i0|i46|i0|qb 0  c=2.98807e-17
c270_3 i0|i46|i0|qb i0|i46|i0|q  c=3.07592e-17
c270_2 i0|i46|i0|qb i0|i44|i0|qb  c=3.55906e-18
c270_1 i0|i46|i0|qb net272  c=6.14999e-18
cg269_3 i0|i46|i0|q 0  c=2.15052e-17
c269_2 i0|i46|i0|q i0|i44|i0|q  c=3.56053e-18
c269_1 i0|i46|i0|q net272  c=1.20485e-17
cg268_3 i0|i44|i3|qb 0  c=2.97054e-17
c268_2 i0|i44|i3|qb i0|i44|i3|q  c=3.0708e-17
c268_1 i0|i44|i3|qb net273  c=5.99196e-18
cg267_2 i0|i44|i3|q 0  c=2.06222e-17
c267_1 i0|i44|i3|q net273  c=1.29959e-17
cg266_3 i0|i44|i2|qb 0  c=3.00508e-17
c266_2 i0|i44|i2|qb i0|i44|i2|q  c=3.06882e-17
c266_1 i0|i44|i2|qb net273  c=5.83386e-18
cg265_2 i0|i44|i2|q 0  c=2.09284e-17
c265_1 i0|i44|i2|q net273  c=1.27096e-17
cg264_3 i0|i44|i1|qb 0  c=2.99377e-17
c264_2 i0|i44|i1|qb i0|i44|i1|q  c=3.07345e-17
c264_1 i0|i44|i1|qb net273  c=5.75256e-18
cg263_2 i0|i44|i1|q 0  c=2.08949e-17
c263_1 i0|i44|i1|q net273  c=1.27792e-17
cg262_3 i0|i44|i0|qb 0  c=3.00613e-17
c262_2 i0|i44|i0|qb i0|i44|i0|q  c=3.06823e-17
c262_1 i0|i44|i0|qb net273  c=5.86113e-18
cg261_2 i0|i44|i0|q 0  c=2.10547e-17
c261_1 i0|i44|i0|q net273  c=1.26447e-17
cg260_4 i0|i38|i3|qb 0  c=2.9637e-17
c260_3 i0|i38|i3|qb i0|i38|i3|q  c=3.07503e-17
c260_2 i0|i38|i3|qb i0|i36|i3|qb  c=3.55906e-18
c260_1 i0|i38|i3|qb net276  c=6.08301e-18
cg259_3 i0|i38|i3|q 0  c=2.09368e-17
c259_2 i0|i38|i3|q i0|i36|i3|q  c=3.56162e-18
c259_1 i0|i38|i3|q net276  c=1.23905e-17
cg258_4 i0|i38|i2|qb 0  c=2.98609e-17
c258_3 i0|i38|i2|qb i0|i38|i2|q  c=3.07667e-17
c258_2 i0|i38|i2|qb i0|i36|i2|qb  c=3.55906e-18
c258_1 i0|i38|i2|qb net276  c=6.10567e-18
cg257_3 i0|i38|i2|q 0  c=2.13814e-17
c257_2 i0|i38|i2|q i0|i36|i2|q  c=3.56053e-18
c257_1 i0|i38|i2|q net276  c=1.20747e-17
cg256_4 i0|i38|i1|qb 0  c=2.98369e-17
c256_3 i0|i38|i1|qb i0|i38|i1|q  c=3.08127e-17
c256_2 i0|i38|i1|qb i0|i36|i1|qb  c=3.55906e-18
c256_1 i0|i38|i1|qb net276  c=6.01587e-18
cg255_3 i0|i38|i1|q 0  c=2.13796e-17
c255_2 i0|i38|i1|q i0|i36|i1|q  c=3.56053e-18
c255_1 i0|i38|i1|q net276  c=1.20928e-17
cg254_4 i0|i38|i0|qb 0  c=2.98947e-17
c254_3 i0|i38|i0|qb i0|i38|i0|q  c=3.07592e-17
c254_2 i0|i38|i0|qb i0|i36|i0|qb  c=3.55906e-18
c254_1 i0|i38|i0|qb net276  c=6.14999e-18
cg253_3 i0|i38|i0|q 0  c=2.14911e-17
c253_2 i0|i38|i0|q i0|i36|i0|q  c=3.56053e-18
c253_1 i0|i38|i0|q net276  c=1.20485e-17
cg252_3 i0|i36|i3|qb 0  c=2.97039e-17
c252_2 i0|i36|i3|qb i0|i36|i3|q  c=3.0708e-17
c252_1 i0|i36|i3|qb net277  c=5.99196e-18
cg251_2 i0|i36|i3|q 0  c=2.06222e-17
c251_1 i0|i36|i3|q net277  c=1.29593e-17
cg250_3 i0|i36|i2|qb 0  c=3.00153e-17
c250_2 i0|i36|i2|qb i0|i36|i2|q  c=3.06805e-17
c250_1 i0|i36|i2|qb net277  c=5.88004e-18
cg249_2 i0|i36|i2|q 0  c=2.09284e-17
c249_1 i0|i36|i2|q net277  c=1.27096e-17
cg248_3 i0|i36|i1|qb 0  c=2.99021e-17
c248_2 i0|i36|i1|qb i0|i36|i1|q  c=3.07268e-17
c248_1 i0|i36|i1|qb net277  c=5.79874e-18
cg247_2 i0|i36|i1|q 0  c=2.08949e-17
c247_1 i0|i36|i1|q net277  c=1.27792e-17
cg246_3 i0|i36|i0|qb 0  c=3.00613e-17
c246_2 i0|i36|i0|qb i0|i36|i0|q  c=3.06823e-17
c246_1 i0|i36|i0|qb net277  c=5.86113e-18
cg245_2 i0|i36|i0|q 0  c=2.10547e-17
c245_1 i0|i36|i0|q net277  c=1.26447e-17
cg244_4 i0|i55|i3|qb 0  c=2.97903e-17
c244_3 i0|i55|i3|qb i0|i55|i3|q  c=3.07484e-17
c244_2 i0|i55|i3|qb i0|i53|i3|qb  c=3.55906e-18
c244_1 i0|i55|i3|qb net264  c=6.16568e-18
cg243_3 i0|i55|i3|q 0  c=2.13819e-17
c243_2 i0|i55|i3|q i0|i53|i3|q  c=3.56053e-18
c243_1 i0|i55|i3|q net264  c=1.20933e-17
cg242_4 i0|i55|i2|qb 0  c=2.98477e-17
c242_3 i0|i55|i2|qb i0|i55|i2|q  c=3.07931e-17
c242_2 i0|i55|i2|qb i0|i53|i2|qb  c=3.55906e-18
c242_1 i0|i55|i2|qb net264  c=6.02086e-18
cg241_3 i0|i55|i2|q 0  c=2.13745e-17
c241_2 i0|i55|i2|q i0|i53|i2|q  c=3.56053e-18
c241_1 i0|i55|i2|q net264  c=1.20954e-17
cg240_4 i0|i55|i1|qb 0  c=2.97968e-17
c240_3 i0|i55|i1|qb i0|i55|i1|q  c=3.07512e-17
c240_2 i0|i55|i1|qb i0|i53|i1|qb  c=3.55906e-18
c240_1 i0|i55|i1|qb net264  c=6.11153e-18
cg239_3 i0|i55|i1|q 0  c=2.14101e-17
c239_2 i0|i55|i1|q i0|i53|i1|q  c=3.56053e-18
c239_1 i0|i55|i1|q net264  c=1.20619e-17
cg238_4 i0|i55|i0|qb 0  c=2.98927e-17
c238_3 i0|i55|i0|qb i0|i55|i0|q  c=3.07306e-17
c238_2 i0|i55|i0|qb i0|i53|i0|qb  c=3.55906e-18
c238_1 i0|i55|i0|qb net264  c=6.06694e-18
cg237_3 i0|i55|i0|q 0  c=2.16835e-17
c237_2 i0|i55|i0|q i0|i53|i0|q  c=3.56053e-18
c237_1 i0|i55|i0|q net264  c=1.20572e-17
cg236_3 i0|i53|i3|qb 0  c=2.9935e-17
c236_2 i0|i53|i3|qb i0|i53|i3|q  c=3.06828e-17
c236_1 i0|i53|i3|qb net269  c=5.89724e-18
cg235_2 i0|i53|i3|q 0  c=2.09048e-17
c235_1 i0|i53|i3|q net269  c=1.27735e-17
cg234_3 i0|i53|i2|qb 0  c=2.98897e-17
c234_2 i0|i53|i2|qb i0|i53|i2|q  c=3.07268e-17
c234_1 i0|i53|i2|qb net269  c=5.82667e-18
cg233_2 i0|i53|i2|q 0  c=2.08971e-17
c233_1 i0|i53|i2|q net269  c=1.27789e-17
cg232_3 i0|i53|i1|qb 0  c=3.00078e-17
c232_2 i0|i53|i1|qb i0|i53|i1|q  c=3.06805e-17
c232_1 i0|i53|i1|qb net269  c=5.87913e-18
cg231_2 i0|i53|i1|q 0  c=2.09445e-17
c231_1 i0|i53|i1|q net269  c=1.26854e-17
cg230_3 i0|i53|i0|qb 0  c=2.99266e-17
c230_2 i0|i53|i0|qb i0|i53|i0|q  c=3.06656e-17
c230_1 i0|i53|i0|qb net269  c=5.79711e-18
cg229_2 i0|i53|i0|q 0  c=2.11355e-17
c229_1 i0|i53|i0|q net269  c=1.27286e-17
cg228_4 i0|i47|i3|qb 0  c=2.97637e-17
c228_3 i0|i47|i3|qb i0|i47|i3|q  c=3.07639e-17
c228_2 i0|i47|i3|qb i0|i45|i3|qb  c=3.55906e-18
c228_1 i0|i47|i3|qb net272  c=6.16568e-18
cg227_3 i0|i47|i3|q 0  c=2.13886e-17
c227_2 i0|i47|i3|q i0|i45|i3|q  c=3.56053e-18
c227_1 i0|i47|i3|q net272  c=1.20933e-17
cg226_4 i0|i47|i2|qb 0  c=2.98212e-17
c226_3 i0|i47|i2|qb i0|i47|i2|q  c=3.08127e-17
c226_2 i0|i47|i2|qb i0|i45|i2|qb  c=3.55906e-18
c226_1 i0|i47|i2|qb net272  c=6.02086e-18
cg225_3 i0|i47|i2|q 0  c=2.1388e-17
c225_2 i0|i47|i2|q i0|i45|i2|q  c=3.56053e-18
c225_1 i0|i47|i2|q net272  c=1.20954e-17
cg224_4 i0|i47|i1|qb 0  c=2.97618e-17
c224_3 i0|i47|i1|qb i0|i47|i1|q  c=3.07645e-17
c224_2 i0|i47|i1|qb i0|i45|i1|qb  c=3.55906e-18
c224_1 i0|i47|i1|qb net272  c=6.11153e-18
cg223_3 i0|i47|i1|q 0  c=2.14113e-17
c223_2 i0|i47|i1|q i0|i45|i1|q  c=3.56053e-18
c223_1 i0|i47|i1|q net272  c=1.20619e-17
cg222_3 i0|i47|i0|qb 0  c=2.98671e-17
c222_2 i0|i47|i0|qb i0|i47|i0|q  c=3.07502e-17
c222_1 i0|i47|i0|qb net272  c=6.06694e-18
cg221_2 i0|i47|i0|q 0  c=2.16824e-17
c221_1 i0|i47|i0|q net272  c=1.20572e-17
cg220_3 i0|i45|i3|qb 0  c=2.99344e-17
c220_2 i0|i45|i3|qb i0|i45|i3|q  c=3.06828e-17
c220_1 i0|i45|i3|qb net273  c=5.89724e-18
cg219_2 i0|i45|i3|q 0  c=2.09061e-17
c219_1 i0|i45|i3|q net273  c=1.27735e-17
cg218_3 i0|i45|i2|qb 0  c=2.99246e-17
c218_2 i0|i45|i2|qb i0|i45|i2|q  c=3.07345e-17
c218_1 i0|i45|i2|qb net273  c=5.78049e-18
cg217_2 i0|i45|i2|q 0  c=2.08984e-17
c217_1 i0|i45|i2|q net273  c=1.27789e-17
cg216_3 i0|i45|i1|qb 0  c=3.00427e-17
c216_2 i0|i45|i1|qb i0|i45|i1|q  c=3.06882e-17
c216_1 i0|i45|i1|qb net273  c=5.83295e-18
cg215_2 i0|i45|i1|q 0  c=2.09458e-17
c215_1 i0|i45|i1|q net273  c=1.26892e-17
cg210_5 i36|i22|i25|net27 0  c=4.05036e-17
c210_4 i36|i22|i25|net27 i36|i22|net54  c=1.1465e-17
c210_3 i36|i22|i25|net27 ln_x5cbbd88253|x5cbbd882345|16  c=3.22429e-18
c210_2 i36|i22|i25|net27 i36|wen  c=2.63329e-17
c210_1 i36|i22|i25|net27 d<3>  c=1.69579e-17
cg209_5 i36|i22|net62 0  c=1.72059e-17
c209_4 i36|i22|net62 ln_x5cbbd88253|x5cbbd882345|17  c=3.37981e-18
c209_3 i36|i22|net62 i36|i22|i24|net27  c=1.60572e-17
c209_2 i36|i22|net62 i36|wen  c=1.68497e-17
c209_1 i36|i22|net62 d<3>  c=1.85698e-17
cg208_4 i36|i22|net54 0  c=2.85682e-17
c208_3 i36|i22|net54 i36|i23|net52  c=1.9694e-18
c208_2 i36|i22|net54 i36|wen  c=2.88819e-18
c208_1 i36|i22|net54 i36|net271  c=1.26009e-17
cg207_5 i36|i22|net52 0  c=2.16364e-17
c207_4 i36|i22|net52 i36|i22|i24|net27  c=2.38159e-17
c207_3 i36|i22|net52 i36|wen  c=4.46621e-18
c207_2 i36|i22|net52 i36|net269  c=1.57528e-17
c207_1 i36|i22|net52 wenb  c=5.50243e-18
cg206_2 ln_x5cbbd88253|x5cbbd882345|17 0  c=2.01957e-18
c206_1 ln_x5cbbd88253|x5cbbd882345|17 i36|i22|i24|net27  c=3.28742e-18
cg205_3 ln_x5cbbd88253|x5cbbd882345|16 0  c=2.00282e-18
c205_2 ln_x5cbbd88253|x5cbbd882345|16 i36|wen  c=3.30963e-18
c205_1 ln_x5cbbd88253|x5cbbd882345|16 d<3>  c=4.31872e-19
cg204_2 i36|i22|i24|net27 0  c=2.82691e-17
c204_1 i36|i22|i24|net27 i36|wen  c=1.88352e-17
cg199_5 i36|i23|i25|net27 0  c=4.04708e-17
c199_4 i36|i23|i25|net27 i36|i23|net54  c=1.14514e-17
c199_3 i36|i23|i25|net27 ln_x5cbbd88253|x5cbbd882344|16  c=3.22429e-18
c199_2 i36|i23|i25|net27 i36|wen  c=2.6277e-17
c199_1 i36|i23|i25|net27 d<2>  c=1.71075e-17
cg198_5 i36|i23|net62 0  c=1.71844e-17
c198_4 i36|i23|net62 ln_x5cbbd88253|x5cbbd882344|17  c=3.37981e-18
c198_3 i36|i23|net62 i36|i23|i24|net27  c=1.60512e-17
c198_2 i36|i23|net62 i36|wen  c=1.68716e-17
c198_1 i36|i23|net62 d<2>  c=1.85819e-17
cg197_4 i36|i23|net54 0  c=2.85603e-17
c197_3 i36|i23|net54 i36|i24|net52  c=1.9691e-18
c197_2 i36|i23|net54 i36|wen  c=2.88817e-18
c197_1 i36|i23|net54 i36|net264  c=1.26099e-17
cg196_4 i36|i23|net52 0  c=2.2591e-17
c196_3 i36|i23|net52 i36|i23|i24|net27  c=2.39901e-17
c196_2 i36|i23|net52 i36|wen  c=3.31088e-18
c196_1 i36|i23|net52 i36|net250  c=1.57907e-17
cg195_2 ln_x5cbbd88253|x5cbbd882344|17 0  c=2.00777e-18
c195_1 ln_x5cbbd88253|x5cbbd882344|17 i36|i23|i24|net27  c=3.28867e-18
cg194_3 ln_x5cbbd88253|x5cbbd882344|16 0  c=2.00282e-18
c194_2 ln_x5cbbd88253|x5cbbd882344|16 i36|wen  c=3.30963e-18
c194_1 ln_x5cbbd88253|x5cbbd882344|16 d<2>  c=4.31872e-19
cg193_2 i36|i23|i24|net27 0  c=2.83517e-17
c193_1 i36|i23|i24|net27 i36|wen  c=1.88445e-17
cg188_5 i36|i24|i25|net27 0  c=4.03723e-17
c188_4 i36|i24|i25|net27 i36|i24|net54  c=1.1435e-17
c188_3 i36|i24|i25|net27 ln_x5cbbd88253|x5cbbd882343|16  c=3.22429e-18
c188_2 i36|i24|i25|net27 i36|wen  c=2.62185e-17
c188_1 i36|i24|i25|net27 d<1>  c=1.7242e-17
cg187_5 i36|i24|net62 0  c=1.71832e-17
c187_4 i36|i24|net62 ln_x5cbbd88253|x5cbbd882343|17  c=3.37981e-18
c187_3 i36|i24|net62 i36|i24|i24|net27  c=1.60794e-17
c187_2 i36|i24|net62 i36|wen  c=1.68716e-17
c187_1 i36|i24|net62 d<1>  c=1.85819e-17
cg186_4 i36|i24|net54 0  c=2.86694e-17
c186_3 i36|i24|net54 i36|i25|net52  c=1.94686e-18
c186_2 i36|i24|net54 i36|wen  c=2.9018e-18
c186_1 i36|i24|net54 i36|net263  c=1.26094e-17
cg185_4 i36|i24|net52 0  c=2.26216e-17
c185_3 i36|i24|net52 i36|i24|i24|net27  c=2.39888e-17
c185_2 i36|i24|net52 i36|wen  c=3.31087e-18
c185_1 i36|i24|net52 i36|net255  c=1.57909e-17
cg184_2 ln_x5cbbd88253|x5cbbd882343|17 0  c=2.01934e-18
c184_1 ln_x5cbbd88253|x5cbbd882343|17 i36|i24|i24|net27  c=3.2916e-18
cg183_3 ln_x5cbbd88253|x5cbbd882343|16 0  c=2.00282e-18
c183_2 ln_x5cbbd88253|x5cbbd882343|16 i36|wen  c=3.30963e-18
c183_1 ln_x5cbbd88253|x5cbbd882343|16 d<1>  c=4.31872e-19
cg182_2 i36|i24|i24|net27 0  c=2.83367e-17
c182_1 i36|i24|i24|net27 i36|wen  c=1.89332e-17
cg177_5 i36|i25|i25|net27 0  c=4.08205e-17
c177_4 i36|i25|i25|net27 i36|i25|net54  c=1.16267e-17
c177_3 i36|i25|i25|net27 ln_x5cbbd88253|x5cbbd882342|16  c=3.22649e-18
c177_2 i36|i25|i25|net27 i36|wen  c=2.43538e-17
c177_1 i36|i25|i25|net27 d<0>  c=1.76223e-17
cg176_5 i36|i25|net62 0  c=1.70962e-17
c176_4 i36|i25|net62 ln_x5cbbd88253|x5cbbd882342|17  c=3.37981e-18
c176_3 i36|i25|net62 i36|i25|i24|net27  c=1.60521e-17
c176_2 i36|i25|net62 i36|wen  c=1.68738e-17
c176_1 i36|i25|net62 d<0>  c=1.86323e-17
cg175_2 i36|i25|net54 0  c=3.36879e-17
c175_1 i36|i25|net54 i36|net262  c=1.26073e-17
cg174_4 i36|i25|net52 0  c=2.27377e-17
c174_3 i36|i25|net52 i36|i25|i24|net27  c=2.3931e-17
c174_2 i36|i25|net52 i36|wen  c=3.34939e-18
c174_1 i36|i25|net52 i36|net254  c=1.58076e-17
cg173_2 ln_x5cbbd88253|x5cbbd882342|17 0  c=2.00591e-18
c173_1 ln_x5cbbd88253|x5cbbd882342|17 i36|i25|i24|net27  c=3.28831e-18
cg172_3 ln_x5cbbd88253|x5cbbd882342|16 0  c=2.00282e-18
c172_2 ln_x5cbbd88253|x5cbbd882342|16 i36|wen  c=3.30963e-18
c172_1 ln_x5cbbd88253|x5cbbd882342|16 d<0>  c=4.82142e-19
cg171_2 i36|i25|i24|net27 0  c=2.83631e-17
c171_1 i36|i25|i24|net27 i36|wen  c=1.88646e-17
cg170_6 i36|wen 0  c=1.9481e-16
c170_5 i36|wen d<0>  c=1.09596e-17
c170_4 i36|wen d<1>  c=1.44288e-17
c170_3 i36|wen d<2>  c=1.42438e-17
c170_2 i36|wen d<3>  c=1.40957e-17
c170_1 i36|wen wenb  c=2.62479e-17
cg169_3 i0|i61|i2|q 0  c=2.19848e-17
c169_2 i0|i61|i2|q i0|i61|i2|qb  c=3.0727e-17
c169_1 i0|i61|i2|q net261  c=1.26551e-17
cg168_3 i0|i61|i1|qb 0  c=3.11028e-17
c168_2 i0|i61|i1|qb i0|i61|i1|q  c=3.06799e-17
c168_1 i0|i61|i1|qb net261  c=5.93597e-18
cg167_2 i0|i61|i1|q 0  c=2.19656e-17
c167_1 i0|i61|i1|q net261  c=1.26844e-17
cg166_3 i0|i61|i0|qb 0  c=3.1068e-17
c166_2 i0|i61|i0|qb i0|i61|i0|q  c=3.06651e-17
c166_1 i0|i61|i0|qb net261  c=5.87545e-18
cg165_2 i0|i61|i0|q 0  c=2.22234e-17
c165_1 i0|i61|i0|q net261  c=1.26598e-17
cg164_3 i0|i60|i3|qb 0  c=3.07896e-17
c164_2 i0|i60|i3|qb i0|i60|i3|q  c=3.07093e-17
c164_1 i0|i60|i3|qb net261  c=6.0432e-18
cg163_2 i0|i60|i3|q 0  c=2.16954e-17
c163_1 i0|i60|i3|q net261  c=1.28449e-17
cg162_3 i0|i60|i2|qb 0  c=3.11847e-17
c162_2 i0|i60|i2|qb i0|i60|i2|q  c=3.06807e-17
c162_1 i0|i60|i2|qb net261  c=5.93381e-18
cg161_2 i0|i60|i2|q 0  c=2.20505e-17
c161_1 i0|i60|i2|q net261  c=1.27457e-17
cg160_3 i0|i60|i1|qb 0  c=3.10005e-17
c160_2 i0|i60|i1|qb i0|i60|i1|q  c=3.07281e-17
c160_1 i0|i60|i1|qb net261  c=5.86033e-18
cg159_2 i0|i60|i1|q 0  c=2.19268e-17
c159_1 i0|i60|i1|q net261  c=1.28451e-17
cg158_3 i0|i60|i0|qb 0  c=3.12006e-17
c158_2 i0|i60|i0|qb i0|i60|i0|q  c=3.06821e-17
c158_1 i0|i60|i0|qb net261  c=5.93943e-18
cg157_2 i0|i60|i0|q 0  c=2.2106e-17
c157_1 i0|i60|i0|q net261  c=1.25524e-17
cg156_3 i0|i31|i3|qb 0  c=3.08649e-17
c156_2 i0|i31|i3|qb i0|i31|i3|q  c=3.06983e-17
c156_1 i0|i31|i3|qb net280  c=6.19535e-18
cg155_2 i0|i31|i3|q 0  c=2.23317e-17
c155_1 i0|i31|i3|q net280  c=1.19351e-17
cg154_3 i0|i31|i2|qb 0  c=3.06277e-17
c154_2 i0|i31|i2|qb i0|i31|i2|q  c=3.07479e-17
c154_1 i0|i31|i2|qb net280  c=6.07541e-18
cg153_2 i0|i31|i2|q 0  c=2.23917e-17
c153_1 i0|i31|i2|q net280  c=1.20414e-17
cg152_3 i0|i31|i1|qb 0  c=3.08255e-17
c152_2 i0|i31|i1|qb i0|i31|i1|q  c=3.07506e-17
c152_1 i0|i31|i1|qb net280  c=6.04383e-18
cg151_2 i0|i31|i1|q 0  c=2.2331e-17
c151_1 i0|i31|i1|q net280  c=1.20322e-17
cg150_3 i0|i31|i0|qb 0  c=3.06526e-17
c150_2 i0|i31|i0|qb i0|i31|i0|q  c=3.06857e-17
c150_1 i0|i31|i0|qb net280  c=6.12244e-18
cg149_2 i0|i31|i0|q 0  c=2.28609e-17
c149_1 i0|i31|i0|q net280  c=1.20665e-17
cg148_3 i0|i30|i3|qb 0  c=3.08024e-17
c148_2 i0|i30|i3|qb i0|i30|i3|q  c=3.07119e-17
c148_1 i0|i30|i3|qb net280  c=6.30814e-18
cg147_2 i0|i30|i3|q 0  c=2.19507e-17
c147_1 i0|i30|i3|q net280  c=1.23579e-17
cg146_3 i0|i30|i2|qb 0  c=3.05752e-17
c146_2 i0|i30|i2|qb i0|i30|i2|q  c=3.07159e-17
c146_1 i0|i30|i2|qb net280  c=6.05629e-18
cg145_3 i0|i30|i2|q 0  c=2.23168e-17
c145_2 i0|i30|i2|q net280  c=1.20186e-17
c145_1 i0|i30|i2|q wenb  c=2.82226e-18
cg144_3 i0|i30|i1|qb 0  c=3.09664e-17
c144_2 i0|i30|i1|qb i0|i30|i1|q  c=3.08127e-17
c144_1 i0|i30|i1|qb net280  c=6.03046e-18
cg143_2 i0|i30|i1|q 0  c=2.23155e-17
c143_1 i0|i30|i1|q net280  c=1.21088e-17
cg142_3 i0|i30|i0|qb 0  c=3.06371e-17
c142_2 i0|i30|i0|qb i0|i30|i0|q  c=3.07038e-17
c142_1 i0|i30|i0|qb net280  c=6.20393e-18
cg141_2 i0|i30|i0|q 0  c=2.24856e-17
c141_1 i0|i30|i0|q net280  c=1.2025e-17
cg140_13 i39|ab<4> 0  c=6.00414e-17
c140_12 i39|ab<4> ln_157  c=1.0868e-17
c140_11 i39|ab<4> ln_155  c=1.01973e-17
c140_10 i39|ab<4> ln_153  c=1.00704e-17
c140_9 i39|ab<4> ln_151  c=1.01465e-17
c140_8 i39|ab<4> net355  c=1.63732e-17
c140_7 i39|ab<4> net225  c=1.48363e-17
c140_6 i39|ab<4> net227  c=1.64258e-17
c140_5 i39|ab<4> net229  c=1.66198e-17
c140_4 i39|ab<4> net280  c=4.53316e-17
c140_3 i39|ab<4> bl<4>  c=4.8878e-17
c140_2 i39|ab<4> wenb  c=1.85643e-17
c140_1 i39|ab<4> a<4>  c=9.33429e-17
cg139_10 i36|ab<4> 0  c=1.65784e-16
c139_9 i36|ab<4> i36|net254  c=2.41115e-17
c139_8 i36|ab<4> i36|net262  c=2.42746e-17
c139_7 i36|ab<4> i36|net255  c=2.3947e-17
c139_6 i36|ab<4> i36|net263  c=2.32813e-17
c139_5 i36|ab<4> i36|net264  c=2.33193e-17
c139_4 i36|ab<4> i36|net250  c=2.4012e-17
c139_3 i36|ab<4> i36|net271  c=2.33315e-17
c139_2 i36|ab<4> i36|net269  c=2.40441e-17
c139_1 i36|ab<4> a<4>  c=1.21519e-16
cg126_2 ln_157 0  c=4.16744e-18
c126_1 ln_157 wenb  c=1.31411e-17
cg125_4 ln_156 0  c=4.01547e-18
c125_3 ln_156 net229  c=8.54715e-19
c125_2 ln_156 wenb  c=9.12875e-18
c125_1 ln_156 a<4>  c=1.40099e-17
cg124_2 ln_155 0  c=4.20899e-18
c124_1 ln_155 wenb  c=1.32759e-17
cg123_4 ln_154 0  c=3.64543e-18
c123_3 ln_154 bl<5>  c=9.15257e-19
c123_2 ln_154 wenb  c=9.07498e-18
c123_1 ln_154 a<4>  c=1.46594e-17
cg122_3 ln_153 0  c=3.37196e-18
c122_2 ln_153 blb<2>  c=7.88897e-19
c122_1 ln_153 wenb  c=1.32962e-17
cg121_4 ln_152 0  c=3.64395e-18
c121_3 ln_152 bl<3>  c=9.15257e-19
c121_2 ln_152 wenb  c=9.07805e-18
c121_1 ln_152 a<4>  c=1.44507e-17
cg120_3 ln_151 0  c=3.41066e-18
c120_2 ln_151 blb<0>  c=7.88897e-19
c120_1 ln_151 wenb  c=1.32759e-17
cg119_4 ln_150 0  c=3.64543e-18
c119_3 ln_150 bl<1>  c=9.15257e-19
c119_2 ln_150 wenb  c=9.07499e-18
c119_1 ln_150 a<4>  c=1.46598e-17
cg118_3 i36|net254 0  c=4.68668e-17
c118_2 i36|net254 bl<0>  c=5.3821e-18
c118_1 i36|net254 a<4>  c=1.4064e-17
cg117_2 i36|net262 0  c=3.60066e-17
c117_1 i36|net262 a<4>  c=9.47407e-18
cg116_3 i36|net255 0  c=4.70457e-17
c116_2 i36|net255 bl<1>  c=5.89828e-18
c116_1 i36|net255 a<4>  c=1.39837e-17
cg115_2 i36|net263 0  c=3.59246e-17
c115_1 i36|net263 a<4>  c=1.1066e-17
cg114_2 i36|net264 0  c=3.64315e-17
c114_1 i36|net264 a<4>  c=1.1109e-17
cg113_3 i36|net250 0  c=4.68925e-17
c113_2 i36|net250 bl<2>  c=6.06097e-18
c113_1 i36|net250 a<4>  c=1.40112e-17
cg112_2 i36|net271 0  c=3.49177e-17
c112_1 i36|net271 a<4>  c=1.12294e-17
cg111_3 i36|net269 0  c=4.54967e-17
c111_2 i36|net269 bl<3>  c=5.25497e-18
c111_1 i36|net269 a<4>  c=1.55161e-17
cg110_15 i11|net699 0  c=1.3705e-16
c110_14 i11|net699 i11|net700  c=5.70099e-17
c110_13 i11|net699 i11|net698  c=3.17653e-17
c110_12 i11|net699 net266  c=1.86988e-17
c110_11 i11|net699 net268  c=1.86657e-17
c110_10 i11|net699 net265  c=1.43584e-17
c110_9 i11|net699 net267  c=1.50509e-17
c110_8 i11|net699 net286  c=1.85269e-17
c110_7 i11|net699 net285  c=1.41982e-17
c110_6 i11|net699 net288  c=1.87205e-17
c110_5 i11|net699 net287  c=1.51289e-17
c110_4 i11|net699 a<3>  c=8.77051e-17
c110_3 i11|net699 a<2>  c=8.40481e-17
c110_2 i11|net699 a<1>  c=3.51411e-17
c110_1 i11|net699 a<0>  c=2.9796e-17
cg109_12 i11|net700 0  c=1.59037e-16
c109_11 i11|net700 net266  c=1.76814e-17
c109_10 i11|net700 net268  c=1.81475e-17
c109_9 i11|net700 net265  c=1.437e-17
c109_8 i11|net700 net267  c=1.55196e-17
c109_7 i11|net700 net282  c=1.81767e-17
c109_6 i11|net700 net284  c=1.81771e-17
c109_5 i11|net700 net281  c=1.5679e-17
c109_4 i11|net700 net283  c=1.56819e-17
c109_3 i11|net700 a<3>  c=6.98372e-17
c109_2 i11|net700 a<2>  c=5.5097e-17
c109_1 i11|net700 a<0>  c=1.97099e-17
cg108_13 i11|net698 0  c=1.5686e-16
c108_12 i11|net698 net266  c=2.48194e-17
c108_11 i11|net698 net265  c=4.46463e-17
c108_10 i11|net698 net282  c=2.47747e-17
c108_9 i11|net698 net286  c=2.47926e-17
c108_8 i11|net698 net281  c=4.3613e-17
c108_7 i11|net698 net285  c=4.37304e-17
c108_6 i11|net698 net290  c=2.50586e-17
c108_5 i11|net698 net289  c=4.40062e-17
c108_4 i11|net698 a<2>  c=3.41535e-17
c108_3 i11|net698 a<1>  c=6.51931e-17
c108_2 i11|net698 a<0>  c=1.57972e-16
c108_1 i11|net698 clk  c=3.57881e-17
cg94_4 i32|i3|net4 0  c=4.47665e-17
c94_3 i32|i3|net4 i32|i2|net4  c=6.84248e-18
c94_2 i32|i3|net4 net265  c=2.19551e-17
c94_1 i32|i3|net4 net261  c=2.4324e-17
cg93_5 i32|i1|net4 0  c=4.08467e-17
c93_4 i32|i1|net4 i32|i2|net4  c=1.02768e-17
c93_3 i32|i1|net4 i32|i0|net4  c=6.79801e-18
c93_2 i32|i1|net4 net267  c=2.18469e-17
c93_1 i32|i1|net4 net263  c=2.42426e-17
cg92_5 i33|i3|net4 0  c=4.07947e-17
c92_4 i33|i3|net4 i32|i0|net4  c=1.02768e-17
c92_3 i33|i3|net4 i33|i2|net4  c=6.79801e-18
c92_2 i33|i3|net4 net281  c=2.18469e-17
c92_1 i33|i3|net4 net269  c=2.42426e-17
cg91_5 i35|i1|net4 0  c=4.05676e-17
c91_4 i35|i1|net4 i35|i0|net4  c=6.92576e-18
c91_3 i35|i1|net4 i35|i2|net4  c=1.02769e-17
c91_2 i35|i1|net4 net291  c=2.18469e-17
c91_1 i35|i1|net4 net279  c=2.42426e-17
cg90_5 i35|i3|net4 0  c=4.07466e-17
c90_4 i35|i3|net4 i35|i2|net4  c=6.86487e-18
c90_3 i35|i3|net4 i34|i0|net4  c=1.02768e-17
c90_2 i35|i3|net4 net289  c=2.18469e-17
c90_1 i35|i3|net4 net277  c=2.42425e-17
cg89_5 i34|i1|net4 0  c=4.08239e-17
c89_4 i34|i1|net4 i34|i0|net4  c=6.79801e-18
c89_3 i34|i1|net4 i34|i2|net4  c=1.02768e-17
c89_2 i34|i1|net4 net287  c=2.18285e-17
c89_1 i34|i1|net4 net275  c=2.42364e-17
cg88_5 i34|i3|net4 0  c=4.07943e-17
c88_4 i34|i3|net4 i34|i2|net4  c=6.79801e-18
c88_3 i34|i3|net4 i33|i0|net4  c=1.02768e-17
c88_2 i34|i3|net4 net285  c=2.18181e-17
c88_1 i34|i3|net4 net273  c=2.42099e-17
cg87_5 i33|i1|net4 0  c=4.0757e-17
c87_4 i33|i1|net4 i33|i2|net4  c=1.02768e-17
c87_3 i33|i1|net4 i33|i0|net4  c=6.79801e-18
c87_2 i33|i1|net4 net283  c=2.18469e-17
c87_1 i33|i1|net4 net271  c=2.42696e-17
cg86_12 i11|net697 0  c=2.16903e-16
c86_11 i11|net697 net265  c=8.6501e-18
c86_10 i11|net697 net267  c=8.24107e-18
c86_9 i11|net697 net281  c=8.40596e-18
c86_8 i11|net697 net283  c=8.67726e-18
c86_7 i11|net697 net285  c=8.28573e-18
c86_6 i11|net697 net287  c=8.27966e-18
c86_5 i11|net697 net289  c=8.40635e-18
c86_4 i11|net697 net291  c=8.74299e-18
c86_3 i11|net697 a<1>  c=2.07292e-17
c86_2 i11|net697 a<0>  c=2.85473e-17
c86_1 i11|net697 clk  c=5.82862e-17
cg85_3 i32|i2|net4 0  c=4.04776e-17
c85_2 i32|i2|net4 net266  c=2.12597e-17
c85_1 i32|i2|net4 net262  c=2.31536e-17
cg84_3 i32|i0|net4 0  c=4.04775e-17
c84_2 i32|i0|net4 net268  c=2.12609e-17
c84_1 i32|i0|net4 net264  c=2.31445e-17
cg83_3 i33|i2|net4 0  c=4.04546e-17
c83_2 i33|i2|net4 net282  c=2.12609e-17
c83_1 i33|i2|net4 net270  c=2.31683e-17
cg82_4 i35|i0|net4 0  c=4.37229e-17
c82_3 i35|i0|net4 net292  c=2.13105e-17
c82_2 i35|i0|net4 net280  c=2.3235e-17
c82_1 i35|i0|net4 a<4>  c=7.09501e-18
cg81_3 i35|i2|net4 0  c=4.04545e-17
c81_2 i35|i2|net4 net290  c=2.12609e-17
c81_1 i35|i2|net4 net278  c=2.31445e-17
cg80_3 i34|i0|net4 0  c=4.04545e-17
c80_2 i34|i0|net4 net288  c=2.12609e-17
c80_1 i34|i0|net4 net276  c=2.31445e-17
cg79_3 i34|i2|net4 0  c=4.04545e-17
c79_2 i34|i2|net4 net286  c=2.12609e-17
c79_1 i34|i2|net4 net274  c=2.31436e-17
cg78_3 i33|i0|net4 0  c=4.04545e-17
c78_2 i33|i0|net4 net284  c=2.12609e-17
c78_1 i33|i0|net4 net272  c=2.31445e-17
cg77_3 i40|i0|net4 0  c=4.69111e-17
c77_2 i40|i0|net4 net229  c=2.18101e-17
c77_1 i40|i0|net4 q<3>  c=2.18549e-17
cg76_3 i40|i1|net4 0  c=4.66937e-17
c76_2 i40|i1|net4 net227  c=2.14943e-17
c76_1 i40|i1|net4 q<2>  c=2.20565e-17
cg75_3 i40|i2|net4 0  c=4.67938e-17
c75_2 i40|i2|net4 net225  c=2.15072e-17
c75_1 i40|i2|net4 q<1>  c=2.19597e-17
cg74_3 i40|i3|net4 0  c=4.62995e-17
c74_2 i40|i3|net4 net355  c=2.15241e-17
c74_1 i40|i3|net4 q<0>  c=2.31862e-17
cg73_3 i0|i61|i3|qb 0  c=3.10279e-17
c73_2 i0|i61|i3|qb i0|i61|i3|q  c=3.06841e-17
c73_1 i0|i61|i3|qb net261  c=5.95092e-18
cg72_2 i0|i61|i3|q 0  c=2.19381e-17
c72_1 i0|i61|i3|q net261  c=1.28409e-17
cg71_2 i0|i61|i2|qb 0  c=3.10246e-17
c71_1 i0|i61|i2|qb net261  c=5.899e-18
cg67_4 net355 0  c=4.82649e-17
c67_3 net355 bl<4>  c=4.35811e-18
c67_2 net355 wenb  c=1.90249e-17
c67_1 net355 a<4>  c=2.14356e-17
cg66_4 net225 0  c=4.96657e-17
c66_3 net225 bl<5>  c=6.50086e-18
c66_2 net225 wenb  c=1.89972e-17
c66_1 net225 a<4>  c=2.26618e-17
cg65_3 net227 0  c=5.12556e-17
c65_2 net227 wenb  c=1.96783e-17
c65_1 net227 a<4>  c=2.14629e-17
cg64_3 net229 0  c=4.32197e-17
c64_2 net229 wenb  c=1.0463e-17
c64_1 net229 a<4>  c=1.91126e-17
cg63_4 net266 0  c=1.05726e-16
c63_3 net266 net265  c=1.49721e-17
c63_2 net266 net267  c=6.34864e-18
c63_1 net266 a<0>  c=9.48759e-18
cg62_5 net268 0  c=1.05445e-16
c62_4 net268 net267  c=1.51767e-17
c62_3 net268 net281  c=6.34996e-18
c62_2 net268 a<1>  c=2.47749e-17
c62_1 net268 a<0>  c=9.45805e-18
cg61_2 net265 0  c=1.08649e-16
c61_1 net265 clk  c=1.28267e-17
cg60_3 net267 0  c=1.0758e-16
c60_2 net267 a<1>  c=4.41814e-17
c60_1 net267 clk  c=1.21336e-17
cg59_5 net282 0  c=1.05903e-16
c59_4 net282 net281  c=1.51817e-17
c59_3 net282 net283  c=6.34996e-18
c59_2 net282 a<2>  c=1.8261e-17
c59_1 net282 a<0>  c=9.46235e-18
cg58_6 net284 0  c=1.0562e-16
c58_5 net284 net283  c=1.51827e-17
c58_4 net284 net285  c=6.35076e-18
c58_3 net284 a<2>  c=1.8564e-17
c58_2 net284 a<1>  c=2.47693e-17
c58_1 net284 a<0>  c=9.45951e-18
cg57_5 net286 0  c=1.04125e-16
c57_4 net286 net285  c=1.55175e-17
c57_3 net286 net287  c=6.37208e-18
c57_2 net286 a<3>  c=1.82747e-17
c57_1 net286 a<0>  c=9.46493e-18
cg56_3 net281 0  c=1.09082e-16
c56_2 net281 a<2>  c=1.38218e-17
c56_1 net281 clk  c=1.28606e-17
cg55_4 net283 0  c=1.07591e-16
c55_3 net283 a<2>  c=1.47649e-17
c55_2 net283 a<1>  c=4.45071e-17
c55_1 net283 clk  c=1.22293e-17
cg54_3 net285 0  c=1.08387e-16
c54_2 net285 a<3>  c=1.43117e-17
c54_1 net285 clk  c=1.26655e-17
cg53_6 net288 0  c=1.03705e-16
c53_5 net288 net287  c=1.56089e-17
c53_4 net288 net289  c=6.37318e-18
c53_3 net288 a<3>  c=1.87487e-17
c53_2 net288 a<1>  c=2.47771e-17
c53_1 net288 a<0>  c=9.46493e-18
cg52_6 net290 0  c=1.02858e-16
c52_5 net290 net289  c=1.56595e-17
c52_4 net290 net291  c=6.37773e-18
c52_3 net290 a<3>  c=1.89378e-17
c52_2 net290 a<2>  c=1.88424e-17
c52_1 net290 a<0>  c=9.46189e-18
cg51_6 net292 0  c=1.03145e-16
c51_5 net292 net291  c=1.5714e-17
c51_4 net292 a<3>  c=1.87404e-17
c51_3 net292 a<2>  c=1.92523e-17
c51_2 net292 a<1>  c=2.51637e-17
c51_1 net292 a<0>  c=9.6089e-18
cg50_4 net287 0  c=1.05216e-16
c50_3 net287 a<3>  c=1.62718e-17
c50_2 net287 a<1>  c=4.4321e-17
c50_1 net287 clk  c=1.24461e-17
cg49_4 net289 0  c=1.05371e-16
c49_3 net289 a<3>  c=1.63724e-17
c49_2 net289 a<2>  c=1.40897e-17
c49_1 net289 clk  c=1.27355e-17
cg48_5 net291 0  c=1.02389e-16
c48_4 net291 a<3>  c=1.64716e-17
c48_3 net291 a<2>  c=1.54047e-17
c48_2 net291 a<1>  c=4.51868e-17
c48_1 net291 clk  c=1.26288e-17
cg47_12 net261 0  c=1.62431e-16
c47_11 net261 blb<1>  c=1.99205e-17
c47_10 net261 blb<2>  c=1.97613e-17
c47_9 net261 blb<3>  c=1.97004e-17
c47_8 net261 blb<4>  c=3.14923e-17
c47_7 net261 blb<5>  c=1.89366e-17
c47_6 net261 bl<6>  c=1.81413e-17
c47_5 net261 blb<6>  c=2.42926e-17
c47_4 net261 blb<7>  c=1.95744e-17
c47_3 net261 bl<0>  c=1.62862e-17
c47_2 net261 blb<0>  c=1.9365e-17
c47_1 net261 bl<2>  c=1.66285e-17
cg46_3 net262 0  c=2.988e-16
c46_2 net262 net263  c=1.1899e-16
c46_1 net262 blb<7>  c=1.88924e-17
cg45_9 net263 0  c=1.74098e-16
c45_8 net263 blb<1>  c=1.98223e-17
c45_7 net263 blb<2>  c=1.84299e-17
c45_6 net263 blb<3>  c=1.94257e-17
c45_5 net263 blb<4>  c=2.02677e-17
c45_4 net263 blb<5>  c=1.88242e-17
c45_3 net263 blb<6>  c=1.98178e-17
c45_2 net263 blb<7>  c=1.93095e-17
c45_1 net263 blb<0>  c=1.87734e-17
cg44_3 net264 0  c=2.99181e-16
c44_2 net264 net269  c=1.18991e-16
c44_1 net264 blb<7>  c=1.88303e-17
cg43_9 net269 0  c=1.7433e-16
c43_8 net269 blb<1>  c=1.98186e-17
c43_7 net269 blb<2>  c=1.84299e-17
c43_6 net269 blb<3>  c=1.94257e-17
c43_5 net269 blb<4>  c=2.02629e-17
c43_4 net269 blb<5>  c=1.88242e-17
c43_3 net269 blb<6>  c=1.98141e-17
c43_2 net269 blb<7>  c=1.93095e-17
c43_1 net269 blb<0>  c=1.87734e-17
cg42_3 net270 0  c=2.99131e-16
c42_2 net270 net271  c=1.18991e-16
c42_1 net270 blb<7>  c=1.88299e-17
cg41_9 net271 0  c=1.7431e-16
c41_8 net271 blb<1>  c=1.98223e-17
c41_7 net271 blb<2>  c=1.84299e-17
c41_6 net271 blb<3>  c=1.94257e-17
c41_5 net271 blb<4>  c=2.02677e-17
c41_4 net271 blb<5>  c=1.88242e-17
c41_3 net271 blb<6>  c=1.98178e-17
c41_2 net271 blb<7>  c=1.93096e-17
c41_1 net271 blb<0>  c=1.87734e-17
cg40_3 net272 0  c=2.99124e-16
c40_2 net272 net273  c=1.18991e-16
c40_1 net272 blb<7>  c=1.88303e-17
cg39_9 net273 0  c=1.74287e-16
c39_8 net273 blb<1>  c=1.98224e-17
c39_7 net273 blb<2>  c=1.84299e-17
c39_6 net273 blb<3>  c=1.94258e-17
c39_5 net273 blb<4>  c=2.02678e-17
c39_4 net273 blb<5>  c=1.88242e-17
c39_3 net273 blb<6>  c=1.98178e-17
c39_2 net273 blb<7>  c=1.93355e-17
c39_1 net273 blb<0>  c=1.87735e-17
cg38_3 net274 0  c=2.991e-16
c38_2 net274 net275  c=1.18991e-16
c38_1 net274 blb<7>  c=1.88741e-17
cg37_9 net275 0  c=1.7433e-16
c37_8 net275 blb<1>  c=1.98223e-17
c37_7 net275 blb<2>  c=1.84299e-17
c37_6 net275 blb<3>  c=1.94257e-17
c37_5 net275 blb<4>  c=2.02677e-17
c37_4 net275 blb<5>  c=1.88242e-17
c37_3 net275 blb<6>  c=1.98178e-17
c37_2 net275 blb<7>  c=1.93599e-17
c37_1 net275 blb<0>  c=1.87734e-17
cg36_3 net276 0  c=2.99074e-16
c36_2 net276 net277  c=1.18991e-16
c36_1 net276 blb<7>  c=1.8874e-17
cg35_9 net277 0  c=1.74173e-16
c35_8 net277 blb<1>  c=1.98223e-17
c35_7 net277 blb<2>  c=1.84299e-17
c35_6 net277 blb<3>  c=1.94257e-17
c35_5 net277 blb<4>  c=2.02677e-17
c35_4 net277 blb<5>  c=1.88242e-17
c35_3 net277 blb<6>  c=1.98178e-17
c35_2 net277 blb<7>  c=1.93649e-17
c35_1 net277 blb<0>  c=1.87734e-17
cg34_3 net278 0  c=2.98916e-16
c34_2 net278 net279  c=1.18957e-16
c34_1 net278 blb<7>  c=1.88826e-17
cg33_9 net279 0  c=1.75926e-16
c33_8 net279 blb<1>  c=1.98169e-17
c33_7 net279 blb<2>  c=1.83938e-17
c33_6 net279 blb<3>  c=1.94257e-17
c33_5 net279 blb<4>  c=2.02276e-17
c33_4 net279 blb<5>  c=1.88242e-17
c33_3 net279 blb<6>  c=1.98124e-17
c33_2 net279 blb<7>  c=1.93633e-17
c33_1 net279 blb<0>  c=1.87373e-17
cg32_7 net280 0  c=2.6166e-16
c32_6 net280 blb<3>  c=1.69062e-17
c32_5 net280 blb<4>  c=1.68326e-17
c32_4 net280 bl<6>  c=1.75692e-17
c32_3 net280 blb<7>  c=1.87124e-17
c32_2 net280 bl<4>  c=1.90558e-17
c32_1 net280 wenb  c=2.04917e-17
cg31_2 q<0> 0  c=1.86685e-17
c31_1 q<0> bl<0>  c=1.60815e-18
cg30_1 d<0> 0  c=3.52419e-17
cg29_2 q<1> 0  c=2.01291e-17
c29_1 q<1> bl<1>  c=3.00567e-18
cg28_1 d<1> 0  c=3.49241e-17
cg27_2 q<2> 0  c=1.89966e-17
c27_1 q<2> bl<3>  c=3.20521e-18
cg26_1 d<2> 0  c=3.46269e-17
cg25_2 q<3> 0  c=2.05559e-17
c25_1 q<3> bl<3>  c=4.02054e-18
cg24_1 d<3> 0  c=3.43175e-17
cg23_4 blb<1> 0  c=3.92416e-16
c23_3 blb<1> bl<1>  c=6.92607e-17
c23_2 blb<1> bl<2>  c=7.63993e-17
c23_1 blb<1> clk  c=3.18637e-17
cg22_5 blb<2> 0  c=3.95221e-16
c22_4 blb<2> blb<4>  c=2.8889e-17
c22_3 blb<2> bl<2>  c=5.35931e-17
c22_2 blb<2> bl<3>  c=1.08324e-16
c22_1 blb<2> clk  c=3.76905e-17
cg21_5 blb<3> 0  c=4.11947e-16
c21_4 blb<3> blb<5>  c=4.34263e-17
c21_3 blb<3> bl<3>  c=5.07524e-17
c21_2 blb<3> bl<4>  c=7.58227e-17
c21_1 blb<3> clk  c=3.29958e-17
cg20_4 blb<4> 0  c=4.36226e-16
c20_3 blb<4> bl<5>  c=7.48889e-17
c20_2 blb<4> bl<4>  c=6.75609e-17
c20_1 blb<4> clk  c=4.75468e-17
cg19_4 blb<5> 0  c=4.06039e-16
c19_3 blb<5> bl<6>  c=8.99465e-17
c19_2 blb<5> bl<5>  c=6.07207e-17
c19_1 blb<5> clk  c=3.62033e-17
cg18_3 bl<6> 0  c=5.04066e-16
c18_2 bl<6> blb<6>  c=5.59627e-17
c18_1 bl<6> clk  c=5.3952e-17
cg17_4 blb<6> 0  c=4.05189e-16
c17_3 blb<6> bl<7>  c=6.77354e-17
c17_2 blb<6> bl<3>  c=3.67413e-17
c17_1 blb<6> clk  c=4.50537e-17
cg16_5 bl<7> 0  c=4.5842e-16
c16_4 bl<7> blb<7>  c=5.69806e-17
c16_3 bl<7> wenb  c=4.25392e-17
c16_2 bl<7> a<4>  c=2.47365e-17
c16_1 bl<7> clk  c=6.48594e-17
cg15_3 blb<7> 0  c=2.68872e-16
c15_2 blb<7> a<4>  c=3.1351e-17
c15_1 blb<7> clk  c=3.40817e-17
cg14_3 bl<0> 0  c=5.61392e-16
c14_2 bl<0> blb<0>  c=6.12806e-17
c14_1 bl<0> clk  c=5.60038e-17
cg13_4 bl<1> 0  c=5.77179e-16
c13_3 bl<1> blb<0>  c=7.39808e-17
c13_2 bl<1> bl<2>  c=2.43154e-17
c13_1 bl<1> clk  c=6.08575e-17
cg12_5 bl<5> 0  c=5.15913e-16
c12_4 bl<5> bl<2>  c=2.53002e-17
c12_3 bl<5> bl<3>  c=3.52565e-17
c12_2 bl<5> a<4>  c=2.62331e-17
c12_1 bl<5> clk  c=6.84875e-17
cg11_2 blb<0> 0  c=3.86402e-16
c11_1 blb<0> clk  c=3.88661e-17
cg10_3 bl<2> 0  c=5.41725e-16
c10_2 bl<2> a<4>  c=5.56272e-17
c10_1 bl<2> clk  c=5.49452e-17
cg9_2 bl<3> 0  c=5.82066e-16
c9_1 bl<3> clk  c=9.71566e-17
cg8_3 bl<4> 0  c=5.43152e-16
c8_2 bl<4> a<4>  c=6.16435e-17
c8_1 bl<4> clk  c=8.17599e-17
cg7_4 a<3> 0  c=2.31538e-16
c7_3 a<3> a<2>  c=7.21775e-17
c7_2 a<3> a<0>  c=2.26126e-17
c7_1 a<3> clk  c=2.88529e-17
cg6_4 a<2> 0  c=1.70722e-16
c6_3 a<2> a<1>  c=4.21104e-17
c6_2 a<2> a<0>  c=6.61466e-17
c6_1 a<2> clk  c=8.50151e-17
cg5_3 a<1> 0  c=1.96717e-16
c5_2 a<1> a<0>  c=3.95745e-17
c5_1 a<1> clk  c=5.90369e-17
cg4_2 a<0> 0  c=1.91777e-16
c4_1 a<0> clk  c=7.91631e-17
cg3_2 wenb 0  c=4.0096e-16
c3_1 wenb a<4>  c=9.31632e-17
cg2_2 a<4> 0  c=3.67099e-16
c2_1 a<4> clk  c=3.32014e-17
cg1_1 clk 0  c=9.06016e-16
.ends top_level

********************************************************************************
* Library          : project_backup
* Cell             : top_level_tb
* View             : schematic
* View Search List : starrc hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
c1 q<1> gnd! c=1f
c3 q<3> gnd! c=1f
c2 q<2> gnd! c=1f
c0 q<0> gnd! c=1f
r33 i_a<4> gnd! r=1meg
rdwenb i_wenb gnd! r=1meg
rdar1 i_a<3> gnd! r=1meg
rdar0 i_a<2> gnd! r=1meg
rdaw1 i_a<1> gnd! r=1meg
rdaw0 i_a<0> gnd! r=1meg
rddw3 i_d<3> gnd! r=1meg
rddw2 i_d<2> gnd! r=1meg
rddw1 i_d<1> gnd! r=1meg
rddw0 i_d<0> gnd! r=1meg
xi34 a<4> i_a<4> inputbuf
xi25 clk net35 inputbuf
xbwenb wenb i_wenb inputbuf
xbar1 a<3> i_a<3> inputbuf
xbar0 a<2> i_a<2> inputbuf
xbaw1 a<1> i_a<1> inputbuf
xbaw0 a<0> i_a<0> inputbuf
xbdw3 d<3> i_d<3> inputbuf
xbdw2 d<2> i_d<2> inputbuf
xbdw1 d<1> i_d<1> inputbuf
xbdw0 d<0> i_d<0> inputbuf
vclk net35 gnd! dc=0 pulse ( 0 'vdd' 0 'clkrise' 'clkrise' '((clkperiod/2)-clkrise)' 'clkperiod'
+  )
vdd vdd! gnd! dc='vdd'
xi35 a<0> a<1> a<2> a<3> a<4> clk d<0> d<1> d<2> d<3> q<0> q<1> q<2> q<3> wenb
+ top_level










.tran 3p '(clkperiod*32)' start=0
.measure tran Qtot INTEG 'i(vdd)' FROM='0' TO='32*clkperiod'
.measure tran Etot PARAM='-Qtot*vdd'
.measure tran EDP PARAM='Etot*clkperiod*32'
.option opfile=1 split_dp=1
.option probe=1
.probe tran v(*) level=1
.probe tran v(a<0>) v(a<1>) v(a<2>) v(a<3>) v(a<4>) v(clk) v(d<0>) v(d<1>)
+ v(d<2>) v(d<3>) v(xi35.bl<0>) v(xi35.bl<1>) v(xi35.bl<2>) v(xi35.bl<3>)
+ v(xi35.bl<4>) v(xi35.bl<5>) v(xi35.bl<6>) v(xi35.bl<7>) v(xi35.blb<0>)
+ v(xi35.blb<1>) v(xi35.blb<2>) v(xi35.blb<3>) v(xi35.blb<4>) v(xi35.blb<5>)
+ v(xi35.blb<6>) v(xi35.blb<7>) v(q<0>) v(q<1>) v(q<2>) v(q<3>) v(wenb)




.end
